-- Internal ROM BIOS
--
-- Set up as a RAM to allow an alternate BIOS to be loaded from
-- and external location, or changed via code.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity romloader is
   port (
      clock_i        : in  std_logic;
      we_n_i         : in  std_logic;
      addr_i         : in  std_logic_vector(14 downto 0);
      data_i         : in  std_logic_vector(7 downto 0);
      data_o         : out std_logic_vector(7 downto 0)
   );
end;

architecture rtl of romloader is

   type ram_t is array(0 to 24575) of std_logic_vector(7 downto 0);
   signal ram_q : ram_t := (
      x"F3", x"ED", x"56", x"C3", x"80", x"00", x"FF", x"FF", -- 0x0000,
      x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0008,
      x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0010,
      x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0018,
      x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0020,
      x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0028,
      x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0030,
      x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0038,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0040,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0048,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0050,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0058,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C3", x"03", -- 0x0060,
      x"01", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0068,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0070,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0078,
      x"31", x"00", x"64", x"CD", x"39", x"12", x"CD", x"45", -- 0x0080,
      x"0F", x"C3", x"00", x"01", x"FF", x"FF", x"FF", x"FF", -- 0x0088,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0090,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0098,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x00F8,
      x"76", x"18", x"FD", x"F5", x"3A", x"06", x"60", x"3C", -- 0x0100,
      x"32", x"06", x"60", x"F1", x"ED", x"45", x"FD", x"21", -- 0x0108,
      x"02", x"00", x"FD", x"39", x"FD", x"7E", x"00", x"D3", -- 0x0110,
      x"BF", x"FD", x"7E", x"01", x"E6", x"3F", x"D3", x"BF", -- 0x0118,
      x"C9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 0x0120,
      x"00", x"3C", x"42", x"A5", x"81", x"A5", x"99", x"42", -- 0x0128,
      x"3C", x"3C", x"7E", x"DB", x"FF", x"FF", x"DB", x"66", -- 0x0130,
      x"3C", x"6C", x"FE", x"FE", x"FE", x"7C", x"38", x"10", -- 0x0138,
      x"00", x"10", x"38", x"7C", x"FE", x"7C", x"38", x"10", -- 0x0140,
      x"00", x"10", x"38", x"54", x"FE", x"54", x"10", x"38", -- 0x0148,
      x"00", x"10", x"38", x"7C", x"FE", x"FE", x"10", x"38", -- 0x0150,
      x"00", x"00", x"00", x"00", x"30", x"30", x"00", x"00", -- 0x0158,
      x"00", x"FF", x"FF", x"FF", x"E7", x"E7", x"FF", x"FF", -- 0x0160,
      x"FF", x"38", x"44", x"82", x"82", x"82", x"44", x"38", -- 0x0168,
      x"00", x"C7", x"BB", x"7D", x"7D", x"7D", x"BB", x"C7", -- 0x0170,
      x"FF", x"0F", x"03", x"05", x"79", x"88", x"88", x"88", -- 0x0178,
      x"70", x"38", x"44", x"44", x"44", x"38", x"10", x"7C", -- 0x0180,
      x"10", x"30", x"28", x"24", x"24", x"28", x"20", x"E0", -- 0x0188,
      x"C0", x"3C", x"24", x"3C", x"24", x"24", x"E4", x"DC", -- 0x0190,
      x"18", x"10", x"54", x"38", x"EE", x"38", x"54", x"10", -- 0x0198,
      x"00", x"10", x"10", x"10", x"7C", x"10", x"10", x"10", -- 0x01A0,
      x"10", x"10", x"10", x"10", x"FF", x"00", x"00", x"00", -- 0x01A8,
      x"00", x"00", x"00", x"00", x"FF", x"10", x"10", x"10", -- 0x01B0,
      x"10", x"10", x"10", x"10", x"F0", x"10", x"10", x"10", -- 0x01B8,
      x"10", x"10", x"10", x"10", x"1F", x"10", x"10", x"10", -- 0x01C0,
      x"10", x"10", x"10", x"10", x"FF", x"10", x"10", x"10", -- 0x01C8,
      x"10", x"10", x"10", x"10", x"10", x"10", x"10", x"10", -- 0x01D0,
      x"10", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", -- 0x01D8,
      x"00", x"00", x"00", x"00", x"1F", x"10", x"10", x"10", -- 0x01E0,
      x"10", x"00", x"00", x"00", x"F0", x"10", x"10", x"10", -- 0x01E8,
      x"10", x"10", x"10", x"10", x"1F", x"00", x"00", x"00", -- 0x01F0,
      x"00", x"10", x"10", x"10", x"F0", x"00", x"00", x"00", -- 0x01F8,
      x"00", x"81", x"42", x"24", x"18", x"18", x"24", x"42", -- 0x0200,
      x"81", x"7E", x"81", x"BD", x"A1", x"A1", x"BD", x"81", -- 0x0208,
      x"7E", x"1F", x"04", x"04", x"04", x"00", x"00", x"00", -- 0x0210,
      x"00", x"44", x"6C", x"54", x"54", x"00", x"00", x"00", -- 0x0218,
      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 0x0220,
      x"00", x"20", x"20", x"20", x"20", x"00", x"00", x"20", -- 0x0228,
      x"00", x"50", x"50", x"50", x"00", x"00", x"00", x"00", -- 0x0230,
      x"00", x"50", x"50", x"F8", x"50", x"F8", x"50", x"50", -- 0x0238,
      x"00", x"20", x"78", x"A0", x"70", x"28", x"F0", x"20", -- 0x0240,
      x"00", x"C0", x"C8", x"10", x"20", x"40", x"98", x"18", -- 0x0248,
      x"00", x"40", x"A0", x"40", x"A8", x"90", x"98", x"60", -- 0x0250,
      x"00", x"10", x"20", x"40", x"00", x"00", x"00", x"00", -- 0x0258,
      x"00", x"10", x"20", x"40", x"40", x"40", x"20", x"10", -- 0x0260,
      x"00", x"40", x"20", x"10", x"10", x"10", x"20", x"40", -- 0x0268,
      x"00", x"20", x"A8", x"70", x"20", x"70", x"A8", x"20", -- 0x0270,
      x"00", x"00", x"20", x"20", x"F8", x"20", x"20", x"00", -- 0x0278,
      x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", -- 0x0280,
      x"40", x"00", x"00", x"00", x"78", x"00", x"00", x"00", -- 0x0288,
      x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"60", -- 0x0290,
      x"00", x"00", x"00", x"08", x"10", x"20", x"40", x"80", -- 0x0298,
      x"00", x"70", x"88", x"98", x"A8", x"C8", x"88", x"70", -- 0x02A0,
      x"00", x"20", x"60", x"A0", x"20", x"20", x"20", x"F0", -- 0x02A8,
      x"00", x"70", x"88", x"08", x"10", x"60", x"80", x"F8", -- 0x02B0,
      x"00", x"70", x"88", x"08", x"30", x"08", x"88", x"70", -- 0x02B8,
      x"00", x"10", x"30", x"50", x"90", x"F8", x"10", x"10", -- 0x02C0,
      x"00", x"F8", x"80", x"E0", x"10", x"08", x"10", x"E0", -- 0x02C8,
      x"00", x"30", x"40", x"80", x"F0", x"88", x"88", x"70", -- 0x02D0,
      x"00", x"F8", x"88", x"10", x"20", x"20", x"20", x"20", -- 0x02D8,
      x"00", x"70", x"88", x"88", x"70", x"88", x"88", x"70", -- 0x02E0,
      x"00", x"70", x"88", x"88", x"78", x"08", x"10", x"60", -- 0x02E8,
      x"00", x"00", x"00", x"20", x"00", x"00", x"20", x"00", -- 0x02F0,
      x"00", x"00", x"00", x"20", x"00", x"00", x"20", x"20", -- 0x02F8,
      x"40", x"18", x"30", x"60", x"C0", x"60", x"30", x"18", -- 0x0300,
      x"00", x"00", x"00", x"F8", x"00", x"F8", x"00", x"00", -- 0x0308,
      x"00", x"C0", x"60", x"30", x"18", x"30", x"60", x"C0", -- 0x0310,
      x"00", x"70", x"88", x"08", x"10", x"20", x"00", x"20", -- 0x0318,
      x"00", x"70", x"88", x"08", x"48", x"A8", x"A8", x"70", -- 0x0320,
      x"00", x"20", x"50", x"88", x"88", x"F8", x"88", x"88", -- 0x0328,
      x"00", x"F0", x"48", x"48", x"70", x"48", x"48", x"F0", -- 0x0330,
      x"00", x"30", x"48", x"80", x"80", x"80", x"48", x"30", -- 0x0338,
      x"00", x"E0", x"50", x"48", x"48", x"48", x"50", x"E0", -- 0x0340,
      x"00", x"F8", x"80", x"80", x"F0", x"80", x"80", x"F8", -- 0x0348,
      x"00", x"F8", x"80", x"80", x"F0", x"80", x"80", x"80", -- 0x0350,
      x"00", x"70", x"88", x"80", x"B8", x"88", x"88", x"70", -- 0x0358,
      x"00", x"88", x"88", x"88", x"F8", x"88", x"88", x"88", -- 0x0360,
      x"00", x"70", x"20", x"20", x"20", x"20", x"20", x"70", -- 0x0368,
      x"00", x"38", x"10", x"10", x"10", x"90", x"90", x"60", -- 0x0370,
      x"00", x"88", x"90", x"A0", x"C0", x"A0", x"90", x"88", -- 0x0378,
      x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"F8", -- 0x0380,
      x"00", x"88", x"D8", x"A8", x"A8", x"88", x"88", x"88", -- 0x0388,
      x"00", x"88", x"C8", x"C8", x"A8", x"98", x"98", x"88", -- 0x0390,
      x"00", x"70", x"88", x"88", x"88", x"88", x"88", x"70", -- 0x0398,
      x"00", x"F0", x"88", x"88", x"F0", x"80", x"80", x"80", -- 0x03A0,
      x"00", x"70", x"88", x"88", x"88", x"A8", x"90", x"68", -- 0x03A8,
      x"00", x"F0", x"88", x"88", x"F0", x"A0", x"90", x"88", -- 0x03B0,
      x"00", x"70", x"88", x"80", x"70", x"08", x"88", x"70", -- 0x03B8,
      x"00", x"F8", x"20", x"20", x"20", x"20", x"20", x"20", -- 0x03C0,
      x"00", x"88", x"88", x"88", x"88", x"88", x"88", x"70", -- 0x03C8,
      x"00", x"88", x"88", x"88", x"88", x"50", x"50", x"20", -- 0x03D0,
      x"00", x"88", x"88", x"88", x"A8", x"A8", x"D8", x"88", -- 0x03D8,
      x"00", x"88", x"88", x"50", x"20", x"50", x"88", x"88", -- 0x03E0,
      x"00", x"88", x"88", x"88", x"70", x"20", x"20", x"20", -- 0x03E8,
      x"00", x"F8", x"08", x"10", x"20", x"40", x"80", x"F8", -- 0x03F0,
      x"00", x"70", x"40", x"40", x"40", x"40", x"40", x"70", -- 0x03F8,
      x"00", x"00", x"00", x"80", x"40", x"20", x"10", x"08", -- 0x0400,
      x"00", x"70", x"10", x"10", x"10", x"10", x"10", x"70", -- 0x0408,
      x"00", x"20", x"50", x"88", x"00", x"00", x"00", x"00", -- 0x0410,
      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F8", -- 0x0418,
      x"00", x"80", x"40", x"20", x"00", x"00", x"00", x"00", -- 0x0420,
      x"00", x"00", x"00", x"70", x"08", x"78", x"88", x"78", -- 0x0428,
      x"00", x"80", x"80", x"B0", x"C8", x"88", x"C8", x"B0", -- 0x0430,
      x"00", x"00", x"00", x"70", x"88", x"80", x"88", x"70", -- 0x0438,
      x"00", x"08", x"08", x"68", x"98", x"88", x"98", x"68", -- 0x0440,
      x"00", x"00", x"00", x"70", x"88", x"F8", x"80", x"70", -- 0x0448,
      x"00", x"10", x"28", x"20", x"F8", x"20", x"20", x"20", -- 0x0450,
      x"00", x"00", x"00", x"68", x"98", x"98", x"68", x"08", -- 0x0458,
      x"70", x"80", x"80", x"F0", x"88", x"88", x"88", x"88", -- 0x0460,
      x"00", x"20", x"00", x"60", x"20", x"20", x"20", x"70", -- 0x0468,
      x"00", x"10", x"00", x"30", x"10", x"10", x"10", x"90", -- 0x0470,
      x"60", x"40", x"40", x"48", x"50", x"60", x"50", x"48", -- 0x0478,
      x"00", x"60", x"20", x"20", x"20", x"20", x"20", x"70", -- 0x0480,
      x"00", x"00", x"00", x"D0", x"A8", x"A8", x"A8", x"A8", -- 0x0488,
      x"00", x"00", x"00", x"B0", x"C8", x"88", x"88", x"88", -- 0x0490,
      x"00", x"00", x"00", x"70", x"88", x"88", x"88", x"70", -- 0x0498,
      x"00", x"00", x"00", x"B0", x"C8", x"C8", x"B0", x"80", -- 0x04A0,
      x"80", x"00", x"00", x"68", x"98", x"98", x"68", x"08", -- 0x04A8,
      x"08", x"00", x"00", x"B0", x"C8", x"80", x"80", x"80", -- 0x04B0,
      x"00", x"00", x"00", x"78", x"80", x"70", x"08", x"F0", -- 0x04B8,
      x"00", x"40", x"40", x"F0", x"40", x"40", x"48", x"30", -- 0x04C0,
      x"00", x"00", x"00", x"90", x"90", x"90", x"90", x"68", -- 0x04C8,
      x"00", x"00", x"00", x"88", x"88", x"88", x"50", x"20", -- 0x04D0,
      x"00", x"00", x"00", x"88", x"A8", x"A8", x"A8", x"50", -- 0x04D8,
      x"00", x"00", x"00", x"88", x"50", x"20", x"50", x"88", -- 0x04E0,
      x"00", x"00", x"00", x"88", x"88", x"98", x"68", x"08", -- 0x04E8,
      x"70", x"00", x"00", x"F8", x"10", x"20", x"40", x"F8", -- 0x04F0,
      x"00", x"18", x"20", x"20", x"40", x"20", x"20", x"18", -- 0x04F8,
      x"00", x"20", x"20", x"20", x"00", x"20", x"20", x"20", -- 0x0500,
      x"00", x"C0", x"20", x"20", x"10", x"20", x"20", x"C0", -- 0x0508,
      x"00", x"40", x"A8", x"10", x"00", x"00", x"00", x"00", -- 0x0510,
      x"00", x"00", x"00", x"20", x"50", x"F8", x"00", x"00", -- 0x0518,
      x"00", x"30", x"48", x"80", x"80", x"80", x"48", x"30", -- 0x0520,
      x"60", x"50", x"00", x"90", x"90", x"90", x"90", x"68", -- 0x0528,
      x"00", x"10", x"20", x"70", x"88", x"F8", x"80", x"70", -- 0x0530,
      x"00", x"20", x"50", x"70", x"08", x"78", x"88", x"78", -- 0x0538,
      x"00", x"10", x"20", x"20", x"50", x"88", x"F8", x"88", -- 0x0540,
      x"00", x"40", x"20", x"70", x"08", x"78", x"88", x"78", -- 0x0548,
      x"00", x"50", x"00", x"00", x"00", x"00", x"00", x"00", -- 0x0550,
      x"00", x"00", x"00", x"70", x"88", x"80", x"88", x"70", -- 0x0558,
      x"20", x"20", x"50", x"70", x"88", x"F8", x"80", x"70", -- 0x0560,
      x"00", x"10", x"20", x"70", x"20", x"20", x"20", x"70", -- 0x0568,
      x"00", x"10", x"20", x"70", x"88", x"88", x"88", x"70", -- 0x0570,
      x"00", x"10", x"20", x"88", x"88", x"88", x"88", x"70", -- 0x0578,
      x"00", x"20", x"50", x"20", x"50", x"88", x"F8", x"88", -- 0x0580,
      x"00", x"01", x"02", x"04", x"08", x"10", x"20", x"40", -- 0x0588,
      x"80", x"80", x"40", x"20", x"10", x"08", x"04", x"02", -- 0x0590,
      x"01", x"00", x"10", x"10", x"FF", x"10", x"10", x"00", -- 0x0598,
      x"00", x"10", x"20", x"F8", x"80", x"F0", x"80", x"F8", -- 0x05A0,
      x"00", x"00", x"00", x"6C", x"12", x"7E", x"90", x"6E", -- 0x05A8,
      x"00", x"3E", x"50", x"90", x"9C", x"F0", x"90", x"9E", -- 0x05B0,
      x"00", x"20", x"50", x"70", x"88", x"88", x"88", x"70", -- 0x05B8,
      x"00", x"50", x"00", x"70", x"88", x"88", x"88", x"70", -- 0x05C0,
      x"00", x"40", x"20", x"70", x"88", x"88", x"88", x"70", -- 0x05C8,
      x"00", x"20", x"50", x"00", x"90", x"90", x"90", x"68", -- 0x05D0,
      x"00", x"40", x"20", x"00", x"90", x"90", x"90", x"68", -- 0x05D8,
      x"00", x"50", x"00", x"88", x"88", x"98", x"68", x"08", -- 0x05E0,
      x"70", x"50", x"00", x"70", x"88", x"88", x"88", x"70", -- 0x05E8,
      x"00", x"50", x"00", x"88", x"88", x"88", x"88", x"70", -- 0x05F0,
      x"00", x"20", x"20", x"78", x"80", x"80", x"78", x"20", -- 0x05F8,
      x"20", x"18", x"24", x"20", x"F8", x"20", x"E2", x"5C", -- 0x0600,
      x"00", x"88", x"50", x"20", x"F8", x"20", x"F8", x"20", -- 0x0608,
      x"00", x"60", x"80", x"9C", x"84", x"88", x"90", x"7C", -- 0x0610,
      x"00", x"18", x"20", x"20", x"F8", x"20", x"20", x"20", -- 0x0618,
      x"40", x"10", x"20", x"70", x"08", x"78", x"88", x"78", -- 0x0620,
      x"00", x"10", x"20", x"00", x"60", x"20", x"20", x"70", -- 0x0628,
      x"00", x"10", x"20", x"70", x"88", x"88", x"88", x"70", -- 0x0630,
      x"00", x"10", x"20", x"90", x"90", x"90", x"90", x"68", -- 0x0638,
      x"00", x"28", x"50", x"B0", x"C8", x"88", x"88", x"88", -- 0x0640,
      x"00", x"28", x"50", x"88", x"C8", x"A8", x"98", x"88", -- 0x0648,
      x"00", x"60", x"90", x"90", x"68", x"00", x"F8", x"00", -- 0x0650,
      x"00", x"60", x"90", x"90", x"60", x"00", x"F0", x"00", -- 0x0658,
      x"00", x"20", x"00", x"20", x"40", x"80", x"88", x"70", -- 0x0660,
      x"00", x"00", x"00", x"00", x"F8", x"80", x"80", x"00", -- 0x0668,
      x"00", x"00", x"00", x"00", x"F8", x"08", x"08", x"00", -- 0x0670,
      x"00", x"84", x"88", x"90", x"A8", x"54", x"84", x"08", -- 0x0678,
      x"1C", x"84", x"88", x"90", x"A8", x"58", x"A8", x"3C", -- 0x0680,
      x"08", x"20", x"00", x"00", x"20", x"20", x"20", x"20", -- 0x0688,
      x"00", x"00", x"12", x"24", x"48", x"90", x"48", x"24", -- 0x0690,
      x"12", x"00", x"90", x"48", x"24", x"12", x"24", x"48", -- 0x0698,
      x"90", x"28", x"50", x"20", x"50", x"88", x"F8", x"88", -- 0x06A0,
      x"00", x"28", x"50", x"70", x"08", x"78", x"88", x"78", -- 0x06A8,
      x"00", x"28", x"50", x"00", x"70", x"20", x"20", x"70", -- 0x06B0,
      x"00", x"28", x"50", x"00", x"20", x"20", x"20", x"70", -- 0x06B8,
      x"00", x"28", x"50", x"70", x"88", x"88", x"88", x"70", -- 0x06C0,
      x"00", x"28", x"50", x"70", x"88", x"88", x"88", x"70", -- 0x06C8,
      x"00", x"28", x"50", x"00", x"88", x"88", x"88", x"70", -- 0x06D0,
      x"00", x"28", x"50", x"00", x"90", x"90", x"90", x"68", -- 0x06D8,
      x"00", x"FC", x"48", x"48", x"48", x"E8", x"08", x"50", -- 0x06E0,
      x"20", x"00", x"A0", x"00", x"A0", x"A0", x"A0", x"20", -- 0x06E8,
      x"40", x"C0", x"44", x"C8", x"54", x"EC", x"54", x"9E", -- 0x06F0,
      x"04", x"10", x"A8", x"40", x"00", x"00", x"00", x"00", -- 0x06F8,
      x"00", x"00", x"20", x"50", x"88", x"50", x"20", x"00", -- 0x0700,
      x"00", x"C4", x"C8", x"10", x"20", x"40", x"B6", x"36", -- 0x0708,
      x"00", x"7C", x"A8", x"A8", x"68", x"28", x"28", x"28", -- 0x0710,
      x"00", x"38", x"40", x"30", x"48", x"48", x"30", x"08", -- 0x0718,
      x"70", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", -- 0x0720,
      x"FF", x"F0", x"F0", x"F0", x"F0", x"0F", x"0F", x"0F", -- 0x0728,
      x"0F", x"00", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0730,
      x"FF", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", -- 0x0738,
      x"00", x"00", x"00", x"00", x"3C", x"3C", x"00", x"00", -- 0x0740,
      x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"00", -- 0x0748,
      x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", -- 0x0750,
      x"C0", x"0F", x"0F", x"0F", x"0F", x"F0", x"F0", x"F0", -- 0x0758,
      x"F0", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", -- 0x0760,
      x"FC", x"03", x"03", x"03", x"03", x"03", x"03", x"03", -- 0x0768,
      x"03", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", x"3F", -- 0x0770,
      x"3F", x"11", x"22", x"44", x"88", x"11", x"22", x"44", -- 0x0778,
      x"88", x"88", x"44", x"22", x"11", x"88", x"44", x"22", -- 0x0780,
      x"11", x"FE", x"7C", x"38", x"10", x"00", x"00", x"00", -- 0x0788,
      x"00", x"00", x"00", x"00", x"00", x"10", x"38", x"7C", -- 0x0790,
      x"FE", x"80", x"C0", x"E0", x"F0", x"E0", x"C0", x"80", -- 0x0798,
      x"00", x"01", x"03", x"07", x"0F", x"07", x"03", x"01", -- 0x07A0,
      x"00", x"FF", x"7E", x"3C", x"18", x"18", x"3C", x"7E", -- 0x07A8,
      x"FF", x"81", x"C3", x"E7", x"FF", x"FF", x"E7", x"C3", -- 0x07B0,
      x"81", x"F0", x"F0", x"F0", x"F0", x"00", x"00", x"00", -- 0x07B8,
      x"00", x"00", x"00", x"00", x"00", x"0F", x"0F", x"0F", -- 0x07C0,
      x"0F", x"0F", x"0F", x"0F", x"0F", x"00", x"00", x"00", -- 0x07C8,
      x"00", x"00", x"00", x"00", x"00", x"F0", x"F0", x"F0", -- 0x07D0,
      x"F0", x"33", x"33", x"CC", x"CC", x"33", x"33", x"CC", -- 0x07D8,
      x"CC", x"00", x"20", x"20", x"50", x"50", x"88", x"F8", -- 0x07E0,
      x"00", x"20", x"20", x"70", x"20", x"70", x"20", x"20", -- 0x07E8,
      x"00", x"00", x"00", x"00", x"50", x"88", x"A8", x"50", -- 0x07F0,
      x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x07F8,
      x"FF", x"00", x"00", x"00", x"00", x"FF", x"FF", x"FF", -- 0x0800,
      x"FF", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", x"F0", -- 0x0808,
      x"F0", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", x"0F", -- 0x0810,
      x"0F", x"FF", x"FF", x"FF", x"FF", x"00", x"00", x"00", -- 0x0818,
      x"00", x"00", x"00", x"68", x"90", x"90", x"90", x"68", -- 0x0820,
      x"00", x"30", x"48", x"48", x"70", x"48", x"48", x"70", -- 0x0828,
      x"C0", x"F8", x"88", x"80", x"80", x"80", x"80", x"80", -- 0x0830,
      x"00", x"F8", x"50", x"50", x"50", x"50", x"50", x"98", -- 0x0838,
      x"00", x"F8", x"88", x"40", x"20", x"40", x"88", x"F8", -- 0x0840,
      x"00", x"00", x"00", x"78", x"90", x"90", x"90", x"60", -- 0x0848,
      x"00", x"00", x"50", x"50", x"50", x"50", x"68", x"80", -- 0x0850,
      x"80", x"00", x"50", x"A0", x"20", x"20", x"20", x"20", -- 0x0858,
      x"00", x"F8", x"20", x"70", x"A8", x"A8", x"70", x"20", -- 0x0860,
      x"F8", x"20", x"50", x"88", x"F8", x"88", x"50", x"20", -- 0x0868,
      x"00", x"70", x"88", x"88", x"88", x"50", x"50", x"D8", -- 0x0870,
      x"00", x"30", x"40", x"40", x"20", x"50", x"50", x"50", -- 0x0878,
      x"20", x"00", x"00", x"00", x"50", x"A8", x"A8", x"50", -- 0x0880,
      x"00", x"08", x"70", x"A8", x"A8", x"A8", x"70", x"80", -- 0x0888,
      x"00", x"38", x"40", x"80", x"F8", x"80", x"40", x"38", -- 0x0890,
      x"00", x"70", x"88", x"88", x"88", x"88", x"88", x"88", -- 0x0898,
      x"00", x"00", x"00", x"F0", x"00", x"F0", x"00", x"F0", -- 0x08A0,
      x"00", x"20", x"20", x"F8", x"20", x"20", x"00", x"F8", -- 0x08A8,
      x"00", x"C0", x"30", x"08", x"30", x"C0", x"00", x"F8", -- 0x08B0,
      x"00", x"18", x"60", x"80", x"60", x"18", x"00", x"F8", -- 0x08B8,
      x"00", x"10", x"28", x"20", x"20", x"20", x"20", x"20", -- 0x08C0,
      x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"A0", -- 0x08C8,
      x"40", x"00", x"20", x"00", x"F8", x"00", x"20", x"00", -- 0x08D0,
      x"00", x"00", x"50", x"A0", x"00", x"50", x"A0", x"00", -- 0x08D8,
      x"00", x"00", x"18", x"24", x"24", x"18", x"00", x"00", -- 0x08E0,
      x"00", x"00", x"30", x"78", x"78", x"30", x"00", x"00", -- 0x08E8,
      x"00", x"00", x"00", x"00", x"00", x"30", x"00", x"00", -- 0x08F0,
      x"00", x"3E", x"20", x"20", x"20", x"A0", x"60", x"20", -- 0x08F8,
      x"00", x"A0", x"50", x"50", x"50", x"00", x"00", x"00", -- 0x0900,
      x"00", x"40", x"A0", x"20", x"40", x"E0", x"00", x"00", -- 0x0908,
      x"00", x"00", x"38", x"38", x"38", x"38", x"38", x"38", -- 0x0910,
      x"00", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0918,
      x"FF", x"30", x"31", x"32", x"33", x"34", x"35", x"36", -- 0x0920,
      x"37", x"38", x"39", x"41", x"42", x"43", x"44", x"45", -- 0x0928,
      x"46", x"00", x"FD", x"21", x"02", x"00", x"FD", x"39", -- 0x0930,
      x"FD", x"7E", x"00", x"D3", x"BF", x"FD", x"7E", x"01", -- 0x0938,
      x"E6", x"3F", x"F6", x"40", x"D3", x"BF", x"C9", x"FD", -- 0x0940,
      x"21", x"03", x"00", x"FD", x"39", x"FD", x"7E", x"00", -- 0x0948,
      x"D3", x"BF", x"FD", x"2B", x"FD", x"7E", x"00", x"E6", -- 0x0950,
      x"3F", x"F6", x"80", x"D3", x"BF", x"C9", x"C1", x"E1", -- 0x0958,
      x"E5", x"C5", x"E5", x"CD", x"32", x"09", x"F1", x"21", -- 0x0960,
      x"04", x"00", x"39", x"56", x"23", x"7E", x"23", x"4E", -- 0x0968,
      x"FE", x"00", x"28", x"01", x"0C", x"47", x"7A", x"D3", -- 0x0970,
      x"BE", x"10", x"FC", x"0D", x"20", x"F9", x"C9", x"C1", -- 0x0978,
      x"E1", x"E5", x"C5", x"E5", x"CD", x"32", x"09", x"F1", -- 0x0980,
      x"21", x"04", x"00", x"39", x"5E", x"23", x"56", x"23", -- 0x0988,
      x"7E", x"23", x"4E", x"FE", x"00", x"28", x"01", x"0C", -- 0x0990,
      x"47", x"79", x"EB", x"0E", x"BE", x"ED", x"B3", x"3D", -- 0x0998,
      x"20", x"FB", x"C9", x"0E", x"00", x"21", x"02", x"00", -- 0x09A0,
      x"39", x"7E", x"23", x"66", x"6F", x"06", x"00", x"09", -- 0x09A8,
      x"7E", x"B7", x"28", x"07", x"79", x"3C", x"28", x"03", -- 0x09B0,
      x"0C", x"18", x"EA", x"69", x"C9", x"C1", x"E1", x"E5", -- 0x09B8,
      x"C5", x"E5", x"CD", x"A3", x"09", x"F1", x"4D", x"59", -- 0x09C0,
      x"16", x"00", x"C5", x"D5", x"21", x"06", x"00", x"39", -- 0x09C8,
      x"4E", x"23", x"46", x"C5", x"2A", x"07", x"60", x"E5", -- 0x09D0,
      x"CD", x"7F", x"09", x"21", x"06", x"00", x"39", x"F9", -- 0x09D8,
      x"C1", x"06", x"00", x"2A", x"07", x"60", x"09", x"22", -- 0x09E0,
      x"07", x"60", x"C9", x"C1", x"E1", x"E5", x"C5", x"E5", -- 0x09E8,
      x"CD", x"BD", x"09", x"F1", x"2A", x"07", x"60", x"23", -- 0x09F0,
      x"22", x"07", x"60", x"2A", x"07", x"60", x"AF", x"BD", -- 0x09F8,
      x"3E", x"03", x"9C", x"30", x"07", x"21", x"00", x"00", -- 0x0A00,
      x"22", x"07", x"60", x"C9", x"3E", x"20", x"D3", x"BE", -- 0x0A08,
      x"C9", x"2A", x"07", x"60", x"01", x"20", x"00", x"09", -- 0x0A10,
      x"22", x"07", x"60", x"AF", x"BD", x"3E", x"03", x"9C", -- 0x0A18,
      x"30", x"07", x"21", x"00", x"00", x"22", x"07", x"60", -- 0x0A20,
      x"C9", x"7D", x"E6", x"E0", x"6F", x"22", x"07", x"60", -- 0x0A28,
      x"C9", x"C1", x"E1", x"E5", x"C5", x"E5", x"CD", x"BD", -- 0x0A30,
      x"09", x"F1", x"C3", x"11", x"0A", x"FD", x"21", x"03", -- 0x0A38,
      x"00", x"FD", x"39", x"FD", x"6E", x"00", x"26", x"00", -- 0x0A40,
      x"29", x"29", x"29", x"29", x"29", x"FD", x"2B", x"FD", -- 0x0A48,
      x"4E", x"00", x"06", x"00", x"09", x"22", x"07", x"60", -- 0x0A50,
      x"C9", x"01", x"21", x"09", x"FD", x"21", x"02", x"00", -- 0x0A58,
      x"FD", x"39", x"FD", x"7E", x"00", x"07", x"07", x"07", -- 0x0A60,
      x"07", x"E6", x"0F", x"E6", x"0F", x"6F", x"26", x"00", -- 0x0A68,
      x"09", x"7E", x"D3", x"BE", x"FD", x"7E", x"00", x"E6", -- 0x0A70,
      x"0F", x"26", x"00", x"6F", x"09", x"7E", x"D3", x"BE", -- 0x0A78,
      x"3E", x"20", x"D3", x"BE", x"C9", x"FD", x"21", x"04", -- 0x0A80,
      x"00", x"FD", x"39", x"FD", x"4E", x"00", x"79", x"F6", -- 0x0A88,
      x"01", x"D3", x"56", x"DB", x"57", x"79", x"D3", x"56", -- 0x0A90,
      x"FD", x"2B", x"FD", x"2B", x"FD", x"7E", x"00", x"D3", -- 0x0A98,
      x"57", x"0E", x"00", x"3E", x"14", x"81", x"5F", x"3E", -- 0x0AA0,
      x"60", x"CE", x"00", x"57", x"1A", x"D3", x"57", x"AF", -- 0x0AA8,
      x"12", x"0C", x"79", x"D6", x"04", x"38", x"EC", x"21", -- 0x0AB0,
      x"03", x"00", x"39", x"7E", x"D3", x"57", x"0E", x"FF", -- 0x0AB8,
      x"DB", x"57", x"47", x"3C", x"20", x"04", x"0D", x"79", -- 0x0AC0,
      x"20", x"F6", x"68", x"C9", x"FD", x"21", x"04", x"00", -- 0x0AC8,
      x"FD", x"39", x"FD", x"7E", x"00", x"F5", x"33", x"FD", -- 0x0AD0,
      x"2B", x"FD", x"7E", x"00", x"F5", x"33", x"FD", x"2B", -- 0x0AD8,
      x"FD", x"7E", x"00", x"F5", x"33", x"CD", x"85", x"0A", -- 0x0AE0,
      x"F1", x"33", x"4D", x"21", x"04", x"00", x"39", x"7E", -- 0x0AE8,
      x"F6", x"01", x"D3", x"56", x"DB", x"57", x"69", x"C9", -- 0x0AF0,
      x"21", x"11", x"60", x"36", x"01", x"21", x"13", x"60", -- 0x0AF8,
      x"36", x"03", x"3E", x"03", x"D3", x"56", x"0E", x"0A", -- 0x0B00,
      x"DB", x"57", x"0D", x"79", x"20", x"FA", x"11", x"95", -- 0x0B08,
      x"02", x"D5", x"3E", x"40", x"F5", x"33", x"CD", x"CC", -- 0x0B10,
      x"0A", x"F1", x"33", x"2D", x"28", x"03", x"2E", x"02", -- 0x0B18,
      x"C9", x"21", x"16", x"60", x"36", x"01", x"21", x"17", -- 0x0B20,
      x"60", x"36", x"AA", x"11", x"87", x"02", x"D5", x"3E", -- 0x0B28,
      x"48", x"F5", x"33", x"CD", x"85", x"0A", x"F1", x"33", -- 0x0B30,
      x"2D", x"20", x"21", x"DB", x"57", x"DB", x"57", x"DB", -- 0x0B38,
      x"57", x"47", x"DB", x"57", x"4F", x"3E", x"03", x"D3", -- 0x0B40,
      x"56", x"DB", x"57", x"10", x"05", x"79", x"D6", x"AA", -- 0x0B48,
      x"28", x"03", x"2E", x"03", x"C9", x"21", x"13", x"60", -- 0x0B50,
      x"36", x"01", x"18", x"43", x"11", x"01", x"02", x"D5", -- 0x0B58,
      x"3E", x"7A", x"F5", x"33", x"CD", x"85", x"0A", x"F1", -- 0x0B60,
      x"33", x"3E", x"01", x"95", x"30", x"09", x"3E", x"03", -- 0x0B68,
      x"D3", x"56", x"DB", x"57", x"2E", x"04", x"C9", x"DB", -- 0x0B70,
      x"57", x"DB", x"57", x"47", x"DB", x"57", x"E6", x"80", -- 0x0B78,
      x"4F", x"04", x"20", x"01", x"0C", x"DB", x"57", x"3E", -- 0x0B80,
      x"03", x"D3", x"56", x"DB", x"57", x"79", x"D6", x"81", -- 0x0B88,
      x"28", x"03", x"2E", x"05", x"C9", x"21", x"11", x"60", -- 0x0B90,
      x"36", x"00", x"21", x"13", x"60", x"36", x"00", x"11", -- 0x0B98,
      x"01", x"02", x"D5", x"3E", x"77", x"F5", x"33", x"CD", -- 0x0BA0,
      x"CC", x"0A", x"F1", x"33", x"45", x"3A", x"11", x"60", -- 0x0BA8,
      x"3D", x"20", x"05", x"21", x"14", x"60", x"36", x"40", -- 0x0BB0,
      x"C5", x"11", x"01", x"02", x"D5", x"3E", x"69", x"F5", -- 0x0BB8,
      x"33", x"CD", x"CC", x"0A", x"F1", x"33", x"7D", x"C1", -- 0x0BC0,
      x"4F", x"3E", x"01", x"B8", x"38", x"03", x"91", x"30", -- 0x0BC8,
      x"1B", x"11", x"01", x"02", x"D5", x"3E", x"41", x"F5", -- 0x0BD0,
      x"33", x"CD", x"CC", x"0A", x"F1", x"33", x"4D", x"3E", -- 0x0BD8,
      x"01", x"91", x"30", x"03", x"2E", x"06", x"C9", x"21", -- 0x0BE0,
      x"13", x"60", x"36", x"02", x"11", x"A8", x"61", x"7A", -- 0x0BE8,
      x"B3", x"28", x"3F", x"79", x"3D", x"20", x"3B", x"3A", -- 0x0BF0,
      x"13", x"60", x"D6", x"02", x"20", x"13", x"D5", x"11", -- 0x0BF8,
      x"01", x"02", x"D5", x"3E", x"41", x"F5", x"33", x"CD", -- 0x0C00,
      x"CC", x"0A", x"F1", x"33", x"7D", x"D1", x"4F", x"18", -- 0x0C08,
      x"1E", x"D5", x"11", x"01", x"02", x"D5", x"3E", x"77", -- 0x0C10,
      x"F5", x"33", x"CD", x"CC", x"0A", x"F1", x"33", x"11", -- 0x0C18,
      x"01", x"02", x"D5", x"3E", x"69", x"F5", x"33", x"CD", -- 0x0C20,
      x"CC", x"0A", x"F1", x"33", x"7D", x"D1", x"4F", x"1B", -- 0x0C28,
      x"18", x"BD", x"7A", x"B3", x"20", x"03", x"2E", x"07", -- 0x0C30,
      x"C9", x"79", x"B7", x"28", x"03", x"2E", x"08", x"C9", -- 0x0C38,
      x"3A", x"11", x"60", x"3D", x"20", x"34", x"11", x"01", -- 0x0C40,
      x"02", x"D5", x"3E", x"7A", x"F5", x"33", x"CD", x"85", -- 0x0C48,
      x"0A", x"F1", x"33", x"3E", x"01", x"95", x"30", x"03", -- 0x0C50,
      x"2E", x"09", x"C9", x"DB", x"57", x"4F", x"DB", x"57", -- 0x0C58,
      x"DB", x"57", x"DB", x"57", x"3E", x"03", x"D3", x"56", -- 0x0C60,
      x"DB", x"57", x"CB", x"71", x"20", x"26", x"21", x"11", -- 0x0C68,
      x"60", x"36", x"00", x"21", x"13", x"60", x"36", x"00", -- 0x0C70,
      x"18", x"1A", x"21", x"16", x"60", x"36", x"02", x"11", -- 0x0C78,
      x"01", x"02", x"D5", x"3E", x"50", x"F5", x"33", x"CD", -- 0x0C80,
      x"CC", x"0A", x"F1", x"33", x"3E", x"01", x"95", x"30", -- 0x0C88,
      x"03", x"2E", x"0A", x"C9", x"2E", x"01", x"C9", x"3A", -- 0x0C90,
      x"11", x"60", x"B7", x"20", x"1A", x"06", x"09", x"FD", -- 0x0C98,
      x"21", x"02", x"00", x"FD", x"39", x"FD", x"CB", x"00", -- 0x0CA0,
      x"26", x"FD", x"CB", x"01", x"16", x"FD", x"CB", x"02", -- 0x0CA8,
      x"16", x"FD", x"CB", x"03", x"16", x"10", x"E8", x"FD", -- 0x0CB0,
      x"21", x"02", x"00", x"FD", x"39", x"FD", x"4E", x"03", -- 0x0CB8,
      x"21", x"14", x"60", x"71", x"23", x"FD", x"4E", x"02", -- 0x0CC0,
      x"71", x"21", x"16", x"60", x"D1", x"C1", x"C5", x"D5", -- 0x0CC8,
      x"70", x"01", x"17", x"60", x"FD", x"7E", x"00", x"02", -- 0x0CD0,
      x"AF", x"57", x"1E", x"01", x"D5", x"3E", x"51", x"F5", -- 0x0CD8,
      x"33", x"CD", x"85", x"0A", x"F1", x"33", x"7D", x"B7", -- 0x0CE0,
      x"28", x"09", x"3E", x"01", x"D3", x"56", x"DB", x"57", -- 0x0CE8,
      x"2E", x"0B", x"C9", x"11", x"A8", x"61", x"DB", x"57", -- 0x0CF0,
      x"47", x"D6", x"FE", x"3E", x"01", x"28", x"01", x"AF", -- 0x0CF8,
      x"4F", x"B7", x"20", x"0A", x"78", x"E6", x"F0", x"28", -- 0x0D00,
      x"05", x"1B", x"7A", x"B3", x"20", x"E8", x"CB", x"41", -- 0x0D08,
      x"20", x"09", x"3E", x"01", x"D3", x"56", x"DB", x"57", -- 0x0D10,
      x"2E", x"0C", x"C9", x"21", x"07", x"00", x"39", x"7E", -- 0x0D18,
      x"2B", x"B6", x"20", x"0E", x"01", x"00", x"02", x"DB", -- 0x0D20,
      x"57", x"D3", x"BE", x"0B", x"78", x"B1", x"20", x"F7", -- 0x0D28,
      x"18", x"13", x"01", x"00", x"02", x"21", x"06", x"00", -- 0x0D30,
      x"39", x"5E", x"23", x"56", x"DB", x"57", x"12", x"0B", -- 0x0D38,
      x"13", x"78", x"B1", x"20", x"F7", x"DB", x"57", x"DB", -- 0x0D40,
      x"57", x"3E", x"01", x"D3", x"56", x"DB", x"57", x"2E", -- 0x0D48,
      x"01", x"C9", x"DB", x"56", x"E6", x"80", x"4F", x"3E", -- 0x0D50,
      x"04", x"FD", x"21", x"00", x"60", x"FD", x"96", x"00", -- 0x0D58,
      x"38", x"76", x"FD", x"5E", x"00", x"16", x"00", x"21", -- 0x0D60,
      x"6D", x"0D", x"19", x"19", x"E9", x"18", x"08", x"18", -- 0x0D68,
      x"36", x"18", x"4F", x"18", x"54", x"18", x"52", x"79", -- 0x0D70,
      x"D6", x"80", x"20", x"24", x"21", x"02", x"00", x"39", -- 0x0D78,
      x"7E", x"B7", x"28", x"54", x"3E", x"14", x"FD", x"21", -- 0x0D80,
      x"01", x"60", x"FD", x"96", x"00", x"30", x"0B", x"FD", -- 0x0D88,
      x"36", x"00", x"00", x"21", x"00", x"60", x"36", x"01", -- 0x0D90,
      x"18", x"3E", x"21", x"01", x"60", x"34", x"18", x"38", -- 0x0D98,
      x"21", x"01", x"60", x"36", x"00", x"18", x"31", x"CD", -- 0x0DA0,
      x"F8", x"0A", x"7D", x"32", x"12", x"60", x"3A", x"12", -- 0x0DA8,
      x"60", x"3D", x"20", x"07", x"21", x"00", x"60", x"36", -- 0x0DB0,
      x"02", x"18", x"1D", x"21", x"00", x"60", x"36", x"03", -- 0x0DB8,
      x"18", x"16", x"21", x"00", x"60", x"36", x"04", x"18", -- 0x0DC0,
      x"0F", x"79", x"D6", x"80", x"28", x"0A", x"21", x"01", -- 0x0DC8,
      x"60", x"36", x"00", x"21", x"00", x"60", x"36", x"00", -- 0x0DD0,
      x"FD", x"21", x"00", x"60", x"FD", x"6E", x"00", x"C9", -- 0x0DD8,
      x"21", x"00", x"80", x"4E", x"23", x"7E", x"FD", x"21", -- 0x0DE0,
      x"02", x"60", x"FD", x"7E", x"00", x"B7", x"28", x"08", -- 0x0DE8,
      x"FD", x"7E", x"00", x"3D", x"28", x"36", x"18", x"47", -- 0x0DF0,
      x"79", x"FE", x"55", x"28", x"04", x"D6", x"AA", x"20", -- 0x0DF8,
      x"24", x"21", x"02", x"00", x"39", x"7E", x"B7", x"28", -- 0x0E00,
      x"36", x"3E", x"28", x"FD", x"21", x"03", x"60", x"FD", -- 0x0E08,
      x"96", x"00", x"30", x"0B", x"FD", x"36", x"00", x"00", -- 0x0E10,
      x"21", x"02", x"60", x"36", x"01", x"18", x"20", x"21", -- 0x0E18,
      x"03", x"60", x"34", x"18", x"1A", x"21", x"03", x"60", -- 0x0E20,
      x"36", x"00", x"18", x"13", x"79", x"FE", x"55", x"28", -- 0x0E28,
      x"0E", x"D6", x"AA", x"28", x"0A", x"21", x"03", x"60", -- 0x0E30,
      x"36", x"00", x"21", x"02", x"60", x"36", x"00", x"FD", -- 0x0E38,
      x"21", x"02", x"60", x"FD", x"6E", x"00", x"C9", x"DB", -- 0x0E40,
      x"FC", x"2F", x"E6", x"4F", x"4F", x"C5", x"21", x"1E", -- 0x0E48,
      x"00", x"E5", x"CD", x"32", x"09", x"F1", x"C1", x"59", -- 0x0E50,
      x"7B", x"E6", x"F0", x"6F", x"26", x"00", x"CB", x"2C", -- 0x0E58,
      x"CB", x"1D", x"CB", x"2C", x"CB", x"1D", x"CB", x"2C", -- 0x0E60,
      x"CB", x"1D", x"CB", x"2C", x"CB", x"1D", x"3E", x"21", -- 0x0E68,
      x"85", x"6F", x"3E", x"09", x"8C", x"67", x"7E", x"D3", -- 0x0E70,
      x"BE", x"7B", x"E6", x"0F", x"5F", x"16", x"00", x"21", -- 0x0E78,
      x"21", x"09", x"19", x"7E", x"D3", x"BE", x"FD", x"21", -- 0x0E80,
      x"04", x"60", x"FD", x"7E", x"00", x"B7", x"28", x"10", -- 0x0E88,
      x"FD", x"7E", x"00", x"3D", x"28", x"39", x"FD", x"7E", -- 0x0E90,
      x"00", x"D6", x"02", x"28", x"6E", x"C3", x"1B", x"0F", -- 0x0E98,
      x"79", x"B7", x"28", x"24", x"21", x"02", x"00", x"39", -- 0x0EA0,
      x"7E", x"B7", x"28", x"74", x"3E", x"04", x"FD", x"21", -- 0x0EA8,
      x"05", x"60", x"FD", x"96", x"00", x"30", x"0B", x"FD", -- 0x0EB0,
      x"36", x"00", x"00", x"21", x"04", x"60", x"36", x"01", -- 0x0EB8,
      x"18", x"5E", x"21", x"05", x"60", x"34", x"18", x"58", -- 0x0EC0,
      x"21", x"05", x"60", x"36", x"00", x"18", x"51", x"21", -- 0x0EC8,
      x"04", x"60", x"36", x"02", x"CB", x"41", x"28", x"07", -- 0x0ED0,
      x"21", x"04", x"60", x"36", x"03", x"18", x"41", x"CB", -- 0x0ED8,
      x"51", x"28", x"07", x"21", x"04", x"60", x"36", x"04", -- 0x0EE0,
      x"18", x"36", x"CB", x"59", x"28", x"07", x"21", x"04", -- 0x0EE8,
      x"60", x"36", x"05", x"18", x"2B", x"CB", x"49", x"28", -- 0x0EF0,
      x"07", x"21", x"04", x"60", x"36", x"06", x"18", x"20", -- 0x0EF8,
      x"CB", x"71", x"28", x"1C", x"21", x"04", x"60", x"36", -- 0x0F00,
      x"07", x"18", x"15", x"79", x"B7", x"20", x"11", x"21", -- 0x0F08,
      x"05", x"60", x"36", x"00", x"21", x"04", x"60", x"36", -- 0x0F10,
      x"00", x"18", x"05", x"21", x"04", x"60", x"36", x"02", -- 0x0F18,
      x"FD", x"21", x"04", x"60", x"FD", x"6E", x"00", x"C9", -- 0x0F20,
      x"11", x"01", x"C0", x"D5", x"CD", x"47", x"09", x"F1", -- 0x0F28,
      x"21", x"3E", x"0F", x"11", x"00", x"60", x"01", x"05", -- 0x0F30,
      x"00", x"ED", x"B0", x"C3", x"00", x"60", x"DB", x"55", -- 0x0F38,
      x"C3", x"00", x"00", x"00", x"C9", x"F5", x"01", x"00", -- 0x0F40,
      x"01", x"C5", x"AF", x"F5", x"33", x"AF", x"F5", x"33", -- 0x0F48,
      x"CD", x"47", x"09", x"F1", x"11", x"01", x"C0", x"D5", -- 0x0F50,
      x"CD", x"47", x"09", x"F1", x"AF", x"57", x"1E", x"02", -- 0x0F58,
      x"D5", x"CD", x"47", x"09", x"F1", x"11", x"03", x"10", -- 0x0F60,
      x"D5", x"CD", x"47", x"09", x"F1", x"11", x"04", x"01", -- 0x0F68,
      x"D5", x"CD", x"47", x"09", x"F1", x"11", x"05", x"0A", -- 0x0F70,
      x"D5", x"CD", x"47", x"09", x"F1", x"11", x"06", x"02", -- 0x0F78,
      x"D5", x"CD", x"47", x"09", x"F1", x"11", x"07", x"1A", -- 0x0F80,
      x"D5", x"CD", x"47", x"09", x"21", x"20", x"00", x"E3", -- 0x0F88,
      x"3E", x"1A", x"F5", x"33", x"21", x"00", x"04", x"E5", -- 0x0F90,
      x"CD", x"5E", x"09", x"F1", x"33", x"21", x"00", x"08", -- 0x0F98,
      x"E3", x"21", x"21", x"01", x"E5", x"21", x"00", x"08", -- 0x0FA0,
      x"E5", x"CD", x"7F", x"09", x"21", x"06", x"00", x"39", -- 0x0FA8,
      x"F9", x"C1", x"3E", x"00", x"D3", x"C0", x"C5", x"21", -- 0x0FB0,
      x"00", x"03", x"E5", x"3E", x"20", x"F5", x"33", x"26", -- 0x0FB8,
      x"00", x"E5", x"CD", x"5E", x"09", x"F1", x"F1", x"33", -- 0x0FC0,
      x"AF", x"F5", x"33", x"AF", x"F5", x"33", x"CD", x"3D", -- 0x0FC8,
      x"0A", x"21", x"BF", x"11", x"E3", x"CD", x"31", x"0A", -- 0x0FD0,
      x"F1", x"11", x"01", x"E0", x"D5", x"CD", x"47", x"09", -- 0x0FD8,
      x"F1", x"C1", x"FD", x"21", x"06", x"60", x"FD", x"7E", -- 0x0FE0,
      x"00", x"91", x"28", x"F6", x"DB", x"BF", x"FD", x"4E", -- 0x0FE8,
      x"00", x"C5", x"11", x"02", x"01", x"D5", x"CD", x"3D", -- 0x0FF0,
      x"0A", x"21", x"D1", x"11", x"E3", x"CD", x"EB", x"09", -- 0x0FF8,
      x"26", x"01", x"E3", x"33", x"CD", x"52", x"0D", x"33", -- 0x1000,
      x"C1", x"FD", x"21", x"01", x"00", x"FD", x"39", x"FD", -- 0x1008,
      x"75", x"00", x"3E", x"04", x"FD", x"96", x"00", x"DA", -- 0x1010,
      x"D1", x"10", x"FD", x"5E", x"00", x"16", x"00", x"21", -- 0x1018,
      x"26", x"10", x"19", x"19", x"19", x"E9", x"C3", x"35", -- 0x1020,
      x"10", x"C3", x"42", x"10", x"C3", x"6A", x"10", x"C3", -- 0x1028,
      x"4F", x"10", x"C3", x"AF", x"10", x"C5", x"21", x"D9", -- 0x1030,
      x"11", x"E5", x"CD", x"BD", x"09", x"F1", x"C1", x"C3", -- 0x1038,
      x"D1", x"10", x"C5", x"21", x"E3", x"11", x"E5", x"CD", -- 0x1040,
      x"BD", x"09", x"F1", x"C1", x"C3", x"D1", x"10", x"C5", -- 0x1048,
      x"21", x"ED", x"11", x"E5", x"CD", x"BD", x"09", x"F1", -- 0x1050,
      x"C1", x"11", x"21", x"09", x"3A", x"12", x"60", x"E6", -- 0x1058,
      x"0F", x"26", x"00", x"6F", x"19", x"7E", x"D3", x"BE", -- 0x1060,
      x"18", x"67", x"C5", x"21", x"F6", x"11", x"E5", x"CD", -- 0x1068,
      x"BD", x"09", x"21", x"A0", x"00", x"E3", x"CD", x"32", -- 0x1070,
      x"09", x"21", x"00", x"64", x"E3", x"21", x"00", x"00", -- 0x1078,
      x"E5", x"21", x"00", x"08", x"E5", x"CD", x"97", x"0C", -- 0x1080,
      x"21", x"06", x"00", x"39", x"F9", x"C1", x"11", x"00", -- 0x1088,
      x"02", x"21", x"00", x"64", x"E3", x"E1", x"E5", x"7E", -- 0x1090,
      x"D3", x"BE", x"1B", x"FD", x"21", x"00", x"00", x"FD", -- 0x1098,
      x"39", x"FD", x"34", x"00", x"20", x"03", x"FD", x"34", -- 0x10A0,
      x"01", x"7A", x"B3", x"20", x"E8", x"18", x"22", x"C5", -- 0x10A8,
      x"21", x"00", x"12", x"E5", x"CD", x"BD", x"09", x"F1", -- 0x10B0,
      x"C1", x"11", x"09", x"60", x"FD", x"21", x"13", x"60", -- 0x10B8,
      x"FD", x"6E", x"00", x"26", x"00", x"29", x"19", x"5E", -- 0x10C0,
      x"23", x"56", x"C5", x"D5", x"CD", x"BD", x"09", x"F1", -- 0x10C8,
      x"C1", x"C5", x"11", x"02", x"02", x"D5", x"CD", x"3D", -- 0x10D0,
      x"0A", x"21", x"06", x"12", x"E3", x"CD", x"EB", x"09", -- 0x10D8,
      x"26", x"01", x"E3", x"33", x"CD", x"E0", x"0D", x"33", -- 0x10E0,
      x"7D", x"C1", x"B7", x"20", x"27", x"C5", x"21", x"0E", -- 0x10E8,
      x"12", x"E5", x"CD", x"BD", x"09", x"21", x"3A", x"00", -- 0x10F0,
      x"E3", x"3E", x"20", x"F5", x"33", x"2A", x"07", x"60", -- 0x10F8,
      x"E5", x"CD", x"5E", x"09", x"F1", x"F1", x"33", x"C1", -- 0x1100,
      x"AF", x"FD", x"21", x"00", x"00", x"FD", x"39", x"FD", -- 0x1108,
      x"77", x"00", x"18", x"20", x"C5", x"21", x"36", x"00", -- 0x1110,
      x"E5", x"21", x"24", x"80", x"E5", x"2A", x"07", x"60", -- 0x1118,
      x"E5", x"CD", x"7F", x"09", x"21", x"06", x"00", x"39", -- 0x1120,
      x"F9", x"C1", x"FD", x"21", x"00", x"00", x"FD", x"39", -- 0x1128,
      x"FD", x"36", x"00", x"01", x"C5", x"3E", x"01", x"F5", -- 0x1130,
      x"33", x"CD", x"47", x"0E", x"33", x"C1", x"FD", x"21", -- 0x1138,
      x"01", x"00", x"FD", x"39", x"FD", x"75", x"00", x"FD", -- 0x1140,
      x"7E", x"00", x"D6", x"03", x"20", x"03", x"05", x"18", -- 0x1148,
      x"0A", x"21", x"01", x"00", x"39", x"7E", x"D6", x"04", -- 0x1150,
      x"20", x"01", x"04", x"3E", x"02", x"90", x"30", x"02", -- 0x1158,
      x"06", x"01", x"78", x"D6", x"01", x"30", x"02", x"06", -- 0x1160,
      x"02", x"C5", x"21", x"20", x"00", x"E5", x"CD", x"32", -- 0x1168,
      x"09", x"F1", x"C1", x"3E", x"20", x"D3", x"BE", x"C5", -- 0x1170,
      x"21", x"40", x"00", x"E5", x"CD", x"32", x"09", x"F1", -- 0x1178,
      x"C1", x"3E", x"20", x"D3", x"BE", x"68", x"26", x"00", -- 0x1180,
      x"29", x"29", x"29", x"29", x"29", x"C5", x"E5", x"CD", -- 0x1188,
      x"32", x"09", x"F1", x"C1", x"3E", x"3E", x"D3", x"BE", -- 0x1190,
      x"FD", x"21", x"01", x"00", x"FD", x"39", x"FD", x"7E", -- 0x1198,
      x"00", x"D6", x"07", x"C2", x"E2", x"0F", x"78", x"D6", -- 0x11A0,
      x"02", x"C2", x"E2", x"0F", x"FD", x"2B", x"FD", x"7E", -- 0x11A8,
      x"00", x"3D", x"C2", x"E2", x"0F", x"C5", x"CD", x"28", -- 0x11B0,
      x"0F", x"C1", x"C3", x"E2", x"0F", x"F1", x"C9", x"44", -- 0x11B8,
      x"65", x"76", x"69", x"63", x"65", x"73", x"20", x"44", -- 0x11C0,
      x"65", x"74", x"65", x"63", x"74", x"65", x"64", x"3A", -- 0x11C8,
      x"00", x"53", x"44", x"43", x"41", x"52", x"44", x"3A", -- 0x11D0,
      x"00", x"4E", x"4F", x"4E", x"45", x"20", x"20", x"20", -- 0x11D8,
      x"20", x"20", x"00", x"49", x"4E", x"49", x"54", x"2E", -- 0x11E0,
      x"2E", x"2E", x"20", x"20", x"00", x"45", x"52", x"52", -- 0x11E8,
      x"4F", x"52", x"3A", x"20", x"20", x"00", x"52", x"45", -- 0x11F0,
      x"41", x"44", x"49", x"4E", x"47", x"2E", x"2E", x"00", -- 0x11F8,
      x"59", x"45", x"53", x"3A", x"20", x"00", x"43", x"41", -- 0x1200,
      x"52", x"54", x"20", x"20", x"3A", x"00", x"4E", x"4F", -- 0x1208,
      x"4E", x"45", x"00", x"53", x"44", x"53", x"43", x"00", -- 0x1210,
      x"53", x"44", x"48", x"43", x"00", x"4D", x"4D", x"43", -- 0x1218,
      x"20", x"00", x"3F", x"3F", x"3F", x"3F", x"00", x"00", -- 0x1220,
      x"00", x"00", x"13", x"12", x"18", x"12", x"1D", x"12", -- 0x1228,
      x"22", x"12", x"01", x"00", x"03", x"00", x"00", x"00", -- 0x1230,
      x"00", x"01", x"12", x"00", x"78", x"B1", x"28", x"08", -- 0x1238,
      x"11", x"06", x"60", x"21", x"27", x"12", x"ED", x"B0", -- 0x1240,
      x"FD", x"21", x"00", x"60", x"FD", x"36", x"00", x"00", -- 0x1248,
      x"FD", x"21", x"01", x"60", x"FD", x"36", x"00", x"00", -- 0x1250,
      x"FD", x"21", x"02", x"60", x"FD", x"36", x"00", x"00", -- 0x1258,
      x"FD", x"21", x"03", x"60", x"FD", x"36", x"00", x"00", -- 0x1260,
      x"FD", x"21", x"04", x"60", x"FD", x"36", x"00", x"00", -- 0x1268,
      x"FD", x"21", x"05", x"60", x"FD", x"36", x"00", x"00", -- 0x1270,
      x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1278,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1280,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1288,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1290,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1298,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x12F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1300,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1308,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1310,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1318,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1320,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1328,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1330,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1338,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1340,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1348,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1350,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1358,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1360,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1368,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1370,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1378,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1380,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1388,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1390,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1398,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x13F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1400,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1408,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1410,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1418,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1420,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1428,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1430,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1438,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1440,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1448,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1450,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1458,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1460,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1468,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1470,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1478,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1480,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1488,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1490,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1498,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x14F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1500,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1508,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1510,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1518,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1520,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1528,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1530,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1538,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1540,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1548,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1550,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1558,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1560,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1568,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1570,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1578,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1580,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1588,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1590,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1598,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x15F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1600,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1608,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1610,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1618,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1620,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1628,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1630,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1638,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1640,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1648,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1650,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1658,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1660,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1668,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1670,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1678,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1680,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1688,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1690,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1698,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x16F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1700,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1708,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1710,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1718,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1720,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1728,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1730,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1738,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1740,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1748,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1750,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1758,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1760,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1768,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1770,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1778,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1780,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1788,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1790,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1798,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x17F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1800,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1808,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1810,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1818,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1820,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1828,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1830,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1838,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1840,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1848,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1850,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1858,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1860,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1868,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1870,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1878,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1880,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1888,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1890,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1898,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x18F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1900,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1908,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1910,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1918,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1920,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1928,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1930,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1938,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1940,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1948,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1950,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1958,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1960,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1968,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1970,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1978,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1980,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1988,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1990,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1998,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x19F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1A98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1AF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1B98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1BF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1C98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1CF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1D98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1DF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1E98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1ED0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1ED8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1EF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1F98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x1FF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2000,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2008,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2010,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2018,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2020,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2028,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2030,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2038,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2040,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2048,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2050,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2058,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2060,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2068,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2070,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2078,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2080,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2088,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2090,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2098,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x20F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2100,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2108,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2110,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2118,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2120,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2128,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2130,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2138,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2140,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2148,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2150,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2158,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2160,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2168,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2170,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2178,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2180,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2188,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2190,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2198,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x21F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2200,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2208,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2210,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2218,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2220,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2228,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2230,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2238,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2240,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2248,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2250,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2258,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2260,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2268,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2270,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2278,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2280,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2288,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2290,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2298,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x22F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2300,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2308,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2310,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2318,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2320,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2328,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2330,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2338,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2340,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2348,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2350,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2358,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2360,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2368,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2370,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2378,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2380,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2388,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2390,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2398,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x23F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2400,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2408,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2410,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2418,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2420,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2428,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2430,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2438,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2440,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2448,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2450,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2458,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2460,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2468,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2470,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2478,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2480,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2488,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2490,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2498,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x24F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2500,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2508,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2510,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2518,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2520,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2528,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2530,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2538,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2540,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2548,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2550,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2558,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2560,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2568,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2570,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2578,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2580,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2588,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2590,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2598,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x25F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2600,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2608,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2610,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2618,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2620,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2628,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2630,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2638,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2640,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2648,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2650,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2658,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2660,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2668,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2670,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2678,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2680,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2688,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2690,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2698,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x26F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2700,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2708,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2710,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2718,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2720,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2728,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2730,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2738,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2740,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2748,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2750,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2758,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2760,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2768,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2770,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2778,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2780,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2788,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2790,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2798,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x27F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2800,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2808,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2810,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2818,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2820,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2828,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2830,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2838,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2840,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2848,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2850,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2858,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2860,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2868,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2870,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2878,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2880,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2888,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2890,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2898,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x28F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2900,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2908,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2910,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2918,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2920,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2928,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2930,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2938,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2940,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2948,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2950,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2958,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2960,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2968,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2970,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2978,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2980,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2988,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2990,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2998,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x29F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2A98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2AF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2B98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2BF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2C98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2CF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2D98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2DF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2E98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2ED0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2ED8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2EF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2F98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x2FF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3000,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3008,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3010,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3018,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3020,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3028,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3030,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3038,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3040,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3048,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3050,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3058,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3060,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3068,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3070,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3078,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3080,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3088,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3090,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3098,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x30F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3100,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3108,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3110,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3118,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3120,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3128,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3130,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3138,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3140,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3148,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3150,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3158,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3160,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3168,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3170,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3178,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3180,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3188,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3190,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3198,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x31F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3200,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3208,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3210,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3218,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3220,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3228,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3230,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3238,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3240,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3248,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3250,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3258,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3260,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3268,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3270,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3278,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3280,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3288,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3290,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3298,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x32F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3300,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3308,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3310,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3318,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3320,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3328,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3330,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3338,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3340,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3348,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3350,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3358,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3360,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3368,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3370,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3378,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3380,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3388,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3390,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3398,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x33F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3400,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3408,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3410,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3418,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3420,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3428,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3430,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3438,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3440,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3448,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3450,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3458,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3460,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3468,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3470,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3478,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3480,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3488,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3490,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3498,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x34F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3500,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3508,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3510,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3518,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3520,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3528,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3530,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3538,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3540,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3548,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3550,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3558,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3560,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3568,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3570,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3578,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3580,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3588,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3590,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3598,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x35F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3600,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3608,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3610,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3618,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3620,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3628,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3630,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3638,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3640,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3648,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3650,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3658,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3660,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3668,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3670,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3678,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3680,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3688,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3690,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3698,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x36F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3700,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3708,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3710,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3718,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3720,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3728,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3730,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3738,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3740,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3748,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3750,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3758,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3760,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3768,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3770,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3778,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3780,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3788,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3790,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3798,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x37F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3800,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3808,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3810,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3818,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3820,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3828,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3830,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3838,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3840,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3848,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3850,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3858,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3860,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3868,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3870,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3878,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3880,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3888,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3890,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3898,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x38F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3900,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3908,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3910,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3918,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3920,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3928,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3930,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3938,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3940,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3948,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3950,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3958,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3960,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3968,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3970,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3978,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3980,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3988,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3990,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3998,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x39F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3A98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3AF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3B98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3BF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3C98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3CF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3D98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3DF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3E98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3ED0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3ED8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3EF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3F98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x3FF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4000,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4008,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4010,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4018,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4020,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4028,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4030,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4038,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4040,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4048,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4050,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4058,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4060,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4068,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4070,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4078,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4080,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4088,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4090,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4098,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x40F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4100,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4108,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4110,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4118,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4120,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4128,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4130,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4138,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4140,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4148,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4150,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4158,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4160,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4168,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4170,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4178,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4180,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4188,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4190,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4198,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x41F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4200,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4208,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4210,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4218,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4220,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4228,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4230,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4238,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4240,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4248,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4250,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4258,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4260,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4268,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4270,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4278,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4280,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4288,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4290,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4298,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x42F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4300,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4308,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4310,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4318,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4320,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4328,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4330,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4338,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4340,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4348,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4350,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4358,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4360,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4368,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4370,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4378,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4380,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4388,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4390,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4398,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x43F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4400,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4408,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4410,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4418,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4420,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4428,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4430,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4438,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4440,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4448,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4450,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4458,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4460,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4468,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4470,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4478,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4480,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4488,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4490,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4498,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x44F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4500,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4508,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4510,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4518,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4520,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4528,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4530,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4538,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4540,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4548,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4550,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4558,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4560,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4568,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4570,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4578,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4580,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4588,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4590,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4598,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x45F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4600,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4608,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4610,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4618,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4620,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4628,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4630,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4638,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4640,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4648,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4650,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4658,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4660,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4668,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4670,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4678,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4680,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4688,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4690,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4698,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x46F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4700,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4708,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4710,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4718,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4720,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4728,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4730,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4738,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4740,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4748,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4750,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4758,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4760,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4768,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4770,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4778,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4780,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4788,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4790,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4798,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x47F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4800,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4808,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4810,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4818,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4820,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4828,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4830,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4838,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4840,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4848,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4850,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4858,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4860,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4868,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4870,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4878,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4880,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4888,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4890,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4898,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x48F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4900,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4908,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4910,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4918,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4920,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4928,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4930,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4938,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4940,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4948,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4950,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4958,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4960,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4968,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4970,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4978,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4980,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4988,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4990,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4998,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x49F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4A98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4AF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4B98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4BF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4C98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4CF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4D98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4DF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4E98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4ED0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4ED8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4EF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4F98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x4FF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5000,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5008,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5010,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5018,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5020,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5028,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5030,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5038,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5040,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5048,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5050,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5058,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5060,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5068,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5070,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5078,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5080,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5088,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5090,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5098,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x50F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5100,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5108,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5110,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5118,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5120,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5128,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5130,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5138,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5140,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5148,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5150,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5158,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5160,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5168,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5170,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5178,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5180,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5188,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5190,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5198,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x51F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5200,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5208,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5210,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5218,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5220,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5228,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5230,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5238,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5240,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5248,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5250,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5258,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5260,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5268,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5270,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5278,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5280,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5288,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5290,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5298,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x52F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5300,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5308,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5310,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5318,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5320,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5328,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5330,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5338,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5340,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5348,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5350,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5358,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5360,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5368,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5370,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5378,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5380,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5388,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5390,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5398,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x53F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5400,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5408,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5410,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5418,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5420,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5428,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5430,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5438,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5440,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5448,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5450,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5458,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5460,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5468,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5470,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5478,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5480,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5488,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5490,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5498,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x54F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5500,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5508,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5510,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5518,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5520,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5528,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5530,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5538,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5540,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5548,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5550,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5558,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5560,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5568,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5570,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5578,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5580,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5588,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5590,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5598,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x55F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5600,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5608,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5610,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5618,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5620,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5628,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5630,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5638,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5640,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5648,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5650,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5658,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5660,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5668,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5670,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5678,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5680,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5688,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5690,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5698,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x56F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5700,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5708,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5710,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5718,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5720,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5728,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5730,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5738,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5740,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5748,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5750,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5758,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5760,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5768,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5770,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5778,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5780,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5788,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5790,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5798,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x57F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5800,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5808,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5810,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5818,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5820,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5828,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5830,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5838,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5840,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5848,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5850,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5858,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5860,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5868,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5870,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5878,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5880,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5888,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5890,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5898,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x58F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5900,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5908,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5910,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5918,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5920,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5928,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5930,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5938,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5940,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5948,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5950,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5958,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5960,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5968,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5970,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5978,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5980,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5988,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5990,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5998,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59A0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59A8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59B0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59B8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59C0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59C8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59D0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59D8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59E0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59E8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59F0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x59F8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5A98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5AF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5B98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5BF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5C98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5CF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5D98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5DF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5E98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5ED0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5ED8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5EF8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F00,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F08,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F10,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F18,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F20,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F28,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F30,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F38,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F40,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F48,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F50,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F58,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F60,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F68,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F70,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F78,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F80,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F88,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F90,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5F98,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FA0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FA8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FB0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FB8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FC0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FC8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"  -- 0x5FF8
   );

begin
   process(clock_i)
   begin
      if rising_edge(clock_i) then
         if we_n_i = '0' then
            ram_q(to_integer(unsigned(addr_i))) <= data_i;
         end if;
         data_o <= ram_q(to_integer(unsigned(addr_i)));
      end if;
   end process;

end rtl;
