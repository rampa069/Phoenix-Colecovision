-- Internal ROM BIOS
--
-- Set up as a RAM to allow an alternate BIOS to be loaded from
-- and external location, or changed via code.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity rombios is
   port (
      clock_i        : in  std_logic;
      we_n_i         : in  std_logic;
      addr_i         : in  std_logic_vector(13 downto 0);
      data_i         : in  std_logic_vector(7 downto 0);
      data_o         : out std_logic_vector(7 downto 0)
   );
end;

architecture rtl of rombios is

   type ram_t is array(0 to 24575) of std_logic_vector(7 downto 0);
   signal ram_q : ram_t := (
      x"31", x"00", x"80", x"C3", x"69", x"00", x"FF", x"FF", -- 0x0000,
      x"C3", x"38", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0008,
      x"C3", x"38", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0010,
      x"C3", x"38", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0018,
      x"C3", x"38", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0020,
      x"C3", x"38", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0028,
      x"C3", x"38", x"00", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0030,
      x"FB", x"ED", x"4D", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0038,
      x"44", x"65", x"61", x"65", x"20", x"4C", x"75", x"6E", -- 0x0040,
      x"61", x"65", x"3A", x"20", x"42", x"65", x"6E", x"65", -- 0x0048,
      x"64", x"69", x"63", x"69", x"74", x"65", x"20", x"6E", -- 0x0050,
      x"6F", x"63", x"74", x"65", x"73", x"20", x"64", x"65", -- 0x0058,
      x"63", x"6F", x"72", x"61", x"2E", x"2E", x"C3", x"90", -- 0x0060,
      x"00", x"21", x"43", x"73", x"36", x"00", x"21", x"00", -- 0x0068,
      x"70", x"11", x"01", x"70", x"01", x"FF", x"1F", x"36", -- 0x0070,
      x"00", x"ED", x"B0", x"31", x"00", x"80", x"CD", x"B0", -- 0x0078,
      x"5F", x"CD", x"61", x"2F", x"CD", x"41", x"0C", x"C7", -- 0x0080,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x0088,
      x"F5", x"E5", x"21", x"43", x"73", x"CB", x"46", x"CA", -- 0x0090,
      x"A8", x"00", x"C5", x"D5", x"FD", x"E5", x"CD", x"27", -- 0x0098,
      x"2F", x"FD", x"E1", x"D1", x"C1", x"C3", x"AA", x"00", -- 0x00A0,
      x"CB", x"FE", x"E1", x"F1", x"ED", x"45", x"DD", x"E5", -- 0x00A8,
      x"DD", x"21", x"04", x"00", x"DD", x"39", x"DD", x"5E", -- 0x00B0,
      x"00", x"DD", x"56", x"01", x"DD", x"6E", x"02", x"DD", -- 0x00B8,
      x"66", x"03", x"DD", x"4E", x"04", x"DD", x"46", x"05", -- 0x00C0,
      x"79", x"B0", x"28", x"02", x"ED", x"B0", x"DD", x"E1", -- 0x00C8,
      x"C9", x"DD", x"E5", x"DD", x"21", x"04", x"00", x"DD", -- 0x00D0,
      x"39", x"DD", x"6E", x"00", x"DD", x"66", x"01", x"DD", -- 0x00D8,
      x"5E", x"02", x"DD", x"4E", x"04", x"DD", x"46", x"05", -- 0x00E0,
      x"79", x"E6", x"03", x"28", x"05", x"73", x"23", x"0B", -- 0x00E8,
      x"18", x"F6", x"78", x"B1", x"28", x"12", x"73", x"23", -- 0x00F0,
      x"73", x"23", x"73", x"23", x"73", x"23", x"79", x"C6", -- 0x00F8,
      x"FC", x"4F", x"78", x"CE", x"FF", x"47", x"18", x"EA", -- 0x0100,
      x"DD", x"E1", x"C9", x"DD", x"E5", x"DD", x"21", x"04", -- 0x0108,
      x"00", x"DD", x"39", x"DD", x"5E", x"00", x"DD", x"56", -- 0x0110,
      x"01", x"DD", x"6E", x"02", x"DD", x"66", x"03", x"DD", -- 0x0118,
      x"4E", x"04", x"DD", x"46", x"05", x"79", x"B0", x"CA", -- 0x0120,
      x"53", x"01", x"7D", x"93", x"7C", x"9A", x"E2", x"33", -- 0x0128,
      x"01", x"EE", x"80", x"F2", x"51", x"01", x"E5", x"79", -- 0x0130,
      x"85", x"6F", x"78", x"8C", x"67", x"7B", x"95", x"7A", -- 0x0138,
      x"9C", x"30", x"0D", x"79", x"83", x"5F", x"78", x"8A", -- 0x0140,
      x"57", x"1B", x"2B", x"ED", x"B8", x"E1", x"18", x"03", -- 0x0148,
      x"E1", x"ED", x"B0", x"DD", x"E1", x"C9", x"3E", x"80", -- 0x0150,
      x"D3", x"BF", x"3E", x"81", x"D3", x"BF", x"3E", x"00", -- 0x0158,
      x"D3", x"BF", x"3E", x"80", x"D3", x"BF", x"3E", x"00", -- 0x0160,
      x"D3", x"BF", x"3E", x"82", x"D3", x"BF", x"3E", x"40", -- 0x0168,
      x"D3", x"BF", x"3E", x"83", x"D3", x"BF", x"3E", x"01", -- 0x0170,
      x"D3", x"BF", x"3E", x"84", x"D3", x"BF", x"3E", x"0E", -- 0x0178,
      x"D3", x"BF", x"3E", x"85", x"D3", x"BF", x"3E", x"03", -- 0x0180,
      x"D3", x"BF", x"3E", x"86", x"D3", x"BF", x"3E", x"E1", -- 0x0188,
      x"D3", x"BF", x"3E", x"87", x"D3", x"BF", x"21", x"46", -- 0x0190,
      x"73", x"36", x"20", x"21", x"02", x"00", x"39", x"7E", -- 0x0198,
      x"F6", x"E0", x"6F", x"C9", x"F0", x"F0", x"F0", x"F0", -- 0x01A0,
      x"F0", x"F0", x"F0", x"F0", x"F0", x"D0", x"80", x"90", -- 0x01A8,
      x"B0", x"30", x"40", x"00", x"1B", x"00", x"38", x"00", -- 0x01B0,
      x"18", x"00", x"00", x"00", x"20", x"DB", x"55", x"31", -- 0x01B8,
      x"B9", x"73", x"2A", x"0A", x"80", x"E9", x"CD", x"13", -- 0x01C0,
      x"3F", x"F5", x"F5", x"DD", x"7E", x"04", x"DD", x"4E", -- 0x01C8,
      x"05", x"D3", x"BF", x"79", x"F6", x"40", x"D3", x"BF", -- 0x01D0,
      x"DD", x"7E", x"06", x"DD", x"86", x"08", x"4F", x"DD", -- 0x01D8,
      x"7E", x"07", x"DD", x"8E", x"09", x"47", x"33", x"33", -- 0x01E0,
      x"C5", x"DD", x"7E", x"06", x"DD", x"96", x"FC", x"DD", -- 0x01E8,
      x"7E", x"07", x"DD", x"9E", x"FD", x"D2", x"75", x"02", -- 0x01F0,
      x"DD", x"6E", x"06", x"DD", x"66", x"07", x"4E", x"23", -- 0x01F8,
      x"DD", x"75", x"06", x"DD", x"74", x"07", x"1E", x"00", -- 0x0200,
      x"79", x"E6", x"C0", x"DD", x"77", x"FE", x"DD", x"36", -- 0x0208,
      x"FF", x"00", x"79", x"E6", x"3F", x"4F", x"0C", x"DD", -- 0x0210,
      x"7E", x"FE", x"B7", x"DD", x"B6", x"FF", x"28", x"26", -- 0x0218,
      x"DD", x"7E", x"FE", x"D6", x"40", x"DD", x"B6", x"FF", -- 0x0220,
      x"28", x"20", x"DD", x"6E", x"06", x"DD", x"66", x"07", -- 0x0228,
      x"DD", x"7E", x"FE", x"D6", x"80", x"DD", x"B6", x"FF", -- 0x0230,
      x"28", x"14", x"DD", x"7E", x"FE", x"D6", x"C0", x"DD", -- 0x0238,
      x"B6", x"FF", x"28", x"14", x"18", x"24", x"1E", x"00", -- 0x0240,
      x"18", x"20", x"1E", x"FF", x"18", x"1C", x"5E", x"23", -- 0x0248,
      x"DD", x"75", x"06", x"DD", x"74", x"07", x"18", x"12", -- 0x0250,
      x"EB", x"79", x"0D", x"B7", x"28", x"8B", x"1A", x"D3", -- 0x0258,
      x"BE", x"13", x"DD", x"73", x"06", x"DD", x"72", x"07", -- 0x0260,
      x"18", x"EF", x"79", x"0D", x"B7", x"CA", x"E9", x"01", -- 0x0268,
      x"7B", x"D3", x"BE", x"18", x"F5", x"DD", x"F9", x"DD", -- 0x0270,
      x"E1", x"C9", x"21", x"43", x"73", x"36", x"00", x"DB", -- 0x0278,
      x"BF", x"32", x"56", x"73", x"21", x"02", x"00", x"39", -- 0x0280,
      x"4E", x"79", x"0D", x"B7", x"C8", x"3A", x"43", x"73", -- 0x0288,
      x"07", x"30", x"FA", x"21", x"43", x"73", x"36", x"00", -- 0x0290,
      x"DB", x"BF", x"32", x"56", x"73", x"18", x"EA", x"CD", -- 0x0298,
      x"13", x"3F", x"21", x"F6", x"FF", x"39", x"F9", x"DD", -- 0x02A0,
      x"36", x"F6", x"FF", x"DD", x"36", x"FB", x"40", x"DD", -- 0x02A8,
      x"36", x"FC", x"01", x"AF", x"DD", x"77", x"FD", x"AF", -- 0x02B0,
      x"DD", x"77", x"FE", x"AF", x"DD", x"77", x"FF", x"3A", -- 0x02B8,
      x"46", x"73", x"D6", x"20", x"20", x"3E", x"21", x"00", -- 0x02C0,
      x"02", x"E5", x"21", x"41", x"64", x"E5", x"21", x"00", -- 0x02C8,
      x"01", x"E5", x"CD", x"2B", x"2E", x"F1", x"F1", x"F1", -- 0x02D0,
      x"21", x"00", x"02", x"E5", x"3E", x"18", x"F5", x"33", -- 0x02D8,
      x"26", x"01", x"E5", x"CD", x"46", x"37", x"F1", x"33", -- 0x02E0,
      x"21", x"C8", x"01", x"E3", x"21", x"C7", x"14", x"E5", -- 0x02E8,
      x"21", x"00", x"09", x"E5", x"CD", x"0A", x"29", x"F1", -- 0x02F0,
      x"F1", x"F1", x"DD", x"36", x"FB", x"00", x"DD", x"36", -- 0x02F8,
      x"FC", x"01", x"18", x"23", x"21", x"68", x"01", x"E5", -- 0x0300,
      x"21", x"41", x"64", x"E5", x"21", x"40", x"01", x"E5", -- 0x0308,
      x"CD", x"2B", x"2E", x"F1", x"F1", x"F1", x"21", x"68", -- 0x0310,
      x"01", x"E5", x"3E", x"20", x"F5", x"33", x"2E", x"40", -- 0x0318,
      x"E5", x"CD", x"46", x"37", x"F1", x"F1", x"33", x"21", -- 0x0320,
      x"46", x"73", x"4E", x"06", x"00", x"03", x"03", x"03", -- 0x0328,
      x"DD", x"7E", x"FB", x"81", x"4F", x"DD", x"7E", x"FC", -- 0x0330,
      x"88", x"47", x"C5", x"21", x"06", x"00", x"E5", x"21", -- 0x0338,
      x"43", x"05", x"E5", x"C5", x"CD", x"0A", x"29", x"F1", -- 0x0340,
      x"F1", x"F1", x"C1", x"FD", x"21", x"46", x"73", x"FD", -- 0x0348,
      x"6E", x"00", x"26", x"00", x"23", x"23", x"09", x"EB", -- 0x0350,
      x"D5", x"21", x"12", x"00", x"E5", x"21", x"4A", x"05", -- 0x0358,
      x"E5", x"D5", x"CD", x"0A", x"29", x"F1", x"F1", x"F1", -- 0x0360,
      x"D1", x"FD", x"21", x"46", x"73", x"FD", x"6E", x"00", -- 0x0368,
      x"26", x"00", x"19", x"EB", x"D5", x"21", x"16", x"00", -- 0x0370,
      x"E5", x"21", x"5D", x"05", x"E5", x"D5", x"CD", x"0A", -- 0x0378,
      x"29", x"F1", x"F1", x"F1", x"D1", x"21", x"12", x"00", -- 0x0380,
      x"19", x"DD", x"75", x"F7", x"DD", x"74", x"F8", x"FD", -- 0x0388,
      x"21", x"46", x"73", x"FD", x"6E", x"00", x"26", x"00", -- 0x0390,
      x"19", x"EB", x"D5", x"21", x"15", x"00", x"E5", x"21", -- 0x0398,
      x"74", x"05", x"E5", x"D5", x"CD", x"0A", x"29", x"F1", -- 0x03A0,
      x"F1", x"F1", x"D1", x"21", x"12", x"00", x"19", x"DD", -- 0x03A8,
      x"75", x"F9", x"DD", x"74", x"FA", x"FD", x"21", x"46", -- 0x03B0,
      x"73", x"FD", x"6E", x"00", x"26", x"00", x"19", x"EB", -- 0x03B8,
      x"D5", x"21", x"0C", x"00", x"E5", x"21", x"8A", x"05", -- 0x03C0,
      x"E5", x"D5", x"CD", x"0A", x"29", x"F1", x"F1", x"F1", -- 0x03C8,
      x"D1", x"FD", x"21", x"46", x"73", x"FD", x"6E", x"00", -- 0x03D0,
      x"26", x"00", x"29", x"19", x"01", x"97", x"05", x"11", -- 0x03D8,
      x"0B", x"00", x"D5", x"C5", x"E5", x"CD", x"0A", x"29", -- 0x03E0,
      x"F1", x"F1", x"F1", x"3E", x"01", x"F5", x"33", x"CD", -- 0x03E8,
      x"7A", x"02", x"33", x"3A", x"45", x"73", x"B7", x"28", -- 0x03F0,
      x"0A", x"DD", x"36", x"FB", x"A3", x"DD", x"36", x"FC", -- 0x03F8,
      x"05", x"18", x"08", x"DD", x"36", x"FB", x"A7", x"DD", -- 0x0400,
      x"36", x"FC", x"05", x"DD", x"4E", x"FB", x"DD", x"46", -- 0x0408,
      x"FC", x"21", x"03", x"00", x"E5", x"C5", x"DD", x"6E", -- 0x0410,
      x"F7", x"DD", x"66", x"F8", x"E5", x"CD", x"0A", x"29", -- 0x0418,
      x"F1", x"F1", x"F1", x"3A", x"44", x"73", x"B7", x"28", -- 0x0420,
      x"05", x"01", x"AB", x"05", x"18", x"03", x"01", x"AE", -- 0x0428,
      x"05", x"21", x"02", x"00", x"E5", x"C5", x"DD", x"6E", -- 0x0430,
      x"F9", x"DD", x"66", x"FA", x"E5", x"CD", x"0A", x"29", -- 0x0438,
      x"F1", x"F1", x"F1", x"DD", x"7E", x"FD", x"B7", x"28", -- 0x0440,
      x"03", x"DD", x"35", x"FD", x"DD", x"7E", x"FE", x"B7", -- 0x0448,
      x"28", x"03", x"DD", x"35", x"FE", x"DD", x"7E", x"FF", -- 0x0450,
      x"B7", x"28", x"03", x"DD", x"35", x"FF", x"CD", x"B1", -- 0x0458,
      x"05", x"FD", x"21", x"39", x"72", x"FD", x"7E", x"00", -- 0x0460,
      x"DD", x"96", x"F6", x"CA", x"EB", x"03", x"FD", x"7E", -- 0x0468,
      x"00", x"DD", x"77", x"F6", x"D6", x"39", x"28", x"78", -- 0x0470,
      x"DD", x"7E", x"F6", x"D6", x"31", x"20", x"23", x"DD", -- 0x0478,
      x"7E", x"FD", x"B7", x"C2", x"EB", x"03", x"FD", x"21", -- 0x0480,
      x"47", x"73", x"FD", x"7E", x"00", x"EE", x"04", x"FD", -- 0x0488,
      x"77", x"00", x"FD", x"7E", x"00", x"D3", x"BF", x"3E", -- 0x0490,
      x"B2", x"D3", x"BF", x"DD", x"36", x"FD", x"0F", x"C3", -- 0x0498,
      x"EB", x"03", x"DD", x"7E", x"F6", x"D6", x"32", x"20", -- 0x04A0,
      x"19", x"DD", x"7E", x"FE", x"B7", x"C2", x"EB", x"03", -- 0x04A8,
      x"3A", x"45", x"73", x"D6", x"01", x"3E", x"00", x"17", -- 0x04B0,
      x"32", x"45", x"73", x"DD", x"36", x"FE", x"0F", x"C3", -- 0x04B8,
      x"EB", x"03", x"DD", x"7E", x"F6", x"D6", x"33", x"20", -- 0x04C0,
      x"19", x"DD", x"7E", x"FF", x"B7", x"C2", x"EB", x"03", -- 0x04C8,
      x"3A", x"44", x"73", x"D6", x"01", x"3E", x"00", x"17", -- 0x04D0,
      x"32", x"44", x"73", x"DD", x"36", x"FF", x"0F", x"C3", -- 0x04D8,
      x"EB", x"03", x"DD", x"7E", x"F6", x"D6", x"30", x"C2", -- 0x04E0,
      x"EB", x"03", x"CD", x"00", x"00", x"C3", x"EB", x"03", -- 0x04E8,
      x"3A", x"46", x"73", x"D6", x"20", x"20", x"35", x"21", -- 0x04F0,
      x"00", x"02", x"E5", x"3E", x"18", x"F5", x"33", x"26", -- 0x04F8,
      x"01", x"E5", x"CD", x"46", x"37", x"F1", x"33", x"21", -- 0x0500,
      x"13", x"05", x"E3", x"21", x"2A", x"0D", x"E5", x"21", -- 0x0508,
      x"00", x"08", x"E5", x"CD", x"C6", x"01", x"F1", x"F1", -- 0x0510,
      x"21", x"00", x"02", x"E3", x"21", x"41", x"64", x"E5", -- 0x0518,
      x"21", x"00", x"01", x"E5", x"CD", x"0A", x"29", x"F1", -- 0x0520,
      x"F1", x"F1", x"18", x"12", x"21", x"68", x"01", x"E5", -- 0x0528,
      x"21", x"41", x"64", x"E5", x"21", x"40", x"01", x"E5", -- 0x0530,
      x"CD", x"0A", x"29", x"F1", x"F1", x"F1", x"DD", x"F9", -- 0x0538,
      x"DD", x"E1", x"C9", x"50", x"52", x"45", x"53", x"53", -- 0x0540,
      x"3A", x"00", x"31", x"20", x"54", x"4F", x"47", x"47", -- 0x0548,
      x"4C", x"45", x"20", x"53", x"43", x"41", x"4E", x"4C", -- 0x0550,
      x"49", x"4E", x"45", x"53", x"00", x"32", x"20", x"54", -- 0x0558,
      x"4F", x"47", x"47", x"4C", x"45", x"20", x"46", x"4C", -- 0x0560,
      x"49", x"43", x"4B", x"45", x"52", x"20", x"28", x"4F", -- 0x0568,
      x"46", x"46", x"29", x"00", x"33", x"20", x"44", x"52", -- 0x0570,
      x"41", x"4D", x"20", x"50", x"41", x"54", x"54", x"45", -- 0x0578,
      x"52", x"4E", x"20", x"28", x"30", x"30", x"30", x"30", -- 0x0580,
      x"29", x"00", x"30", x"20", x"53", x"4F", x"46", x"54", -- 0x0588,
      x"20", x"52", x"45", x"53", x"45", x"54", x"00", x"39", -- 0x0590,
      x"20", x"45", x"58", x"49", x"54", x"20", x"4D", x"45", -- 0x0598,
      x"4E", x"55", x"00", x"4F", x"4E", x"20", x"00", x"4F", -- 0x05A0,
      x"46", x"46", x"00", x"46", x"46", x"00", x"30", x"30", -- 0x05A8,
      x"00", x"3E", x"01", x"F5", x"33", x"CD", x"4B", x"29", -- 0x05B0,
      x"33", x"3A", x"39", x"72", x"3C", x"20", x"14", x"3A", -- 0x05B8,
      x"3B", x"72", x"B7", x"20", x"0E", x"3A", x"3A", x"72", -- 0x05C0,
      x"B7", x"20", x"08", x"3E", x"02", x"F5", x"33", x"CD", -- 0x05C8,
      x"4B", x"29", x"33", x"3A", x"C2", x"66", x"B7", x"C0", -- 0x05D0,
      x"3A", x"C1", x"66", x"FD", x"21", x"39", x"72", x"FD", -- 0x05D8,
      x"96", x"00", x"C8", x"FD", x"7E", x"00", x"FD", x"21", -- 0x05E0,
      x"C1", x"66", x"FD", x"77", x"00", x"FD", x"21", x"39", -- 0x05E8,
      x"72", x"FD", x"7E", x"00", x"D6", x"2A", x"28", x"07", -- 0x05F0,
      x"FD", x"7E", x"00", x"D6", x"23", x"20", x"0E", x"21", -- 0x05F8,
      x"C2", x"66", x"36", x"01", x"CD", x"9F", x"02", x"21", -- 0x0600,
      x"C2", x"66", x"36", x"00", x"C9", x"FD", x"21", x"39", -- 0x0608,
      x"72", x"FD", x"7E", x"00", x"D6", x"30", x"CA", x"47", -- 0x0610,
      x"24", x"18", x"03", x"C3", x"47", x"24", x"3A", x"39", -- 0x0618,
      x"72", x"D6", x"31", x"C0", x"3A", x"4F", x"73", x"D6", -- 0x0620,
      x"01", x"3E", x"00", x"17", x"32", x"4F", x"73", x"21", -- 0x0628,
      x"3B", x"72", x"36", x"80", x"C9", x"CD", x"13", x"3F", -- 0x0630,
      x"F5", x"DD", x"4E", x"06", x"DD", x"46", x"07", x"DD", -- 0x0638,
      x"5E", x"04", x"DD", x"56", x"05", x"0A", x"B7", x"28", -- 0x0640,
      x"2F", x"03", x"C6", x"E3", x"6F", x"26", x"00", x"29", -- 0x0648,
      x"29", x"29", x"D5", x"11", x"AF", x"14", x"19", x"D1", -- 0x0650,
      x"33", x"33", x"E5", x"C5", x"D5", x"21", x"08", x"00", -- 0x0658,
      x"E5", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"E5", -- 0x0660,
      x"D5", x"CD", x"0A", x"29", x"F1", x"F1", x"F1", x"D1", -- 0x0668,
      x"C1", x"21", x"10", x"00", x"19", x"EB", x"18", x"CD", -- 0x0670,
      x"F1", x"DD", x"E1", x"C9", x"CD", x"13", x"3F", x"21", -- 0x0678,
      x"F1", x"FF", x"39", x"F9", x"DD", x"36", x"F1", x"01", -- 0x0680,
      x"DD", x"7E", x"04", x"DD", x"77", x"FD", x"DD", x"7E", -- 0x0688,
      x"05", x"DD", x"77", x"FE", x"DD", x"5E", x"06", x"DD", -- 0x0690,
      x"56", x"07", x"1A", x"B7", x"CA", x"76", x"07", x"DD", -- 0x0698,
      x"7E", x"FD", x"D3", x"BF", x"DD", x"7E", x"FE", x"F6", -- 0x06A0,
      x"40", x"D3", x"BF", x"DD", x"73", x"F2", x"DD", x"72", -- 0x06A8,
      x"F3", x"21", x"01", x"00", x"19", x"DD", x"75", x"F4", -- 0x06B0,
      x"DD", x"74", x"F5", x"DD", x"7E", x"F4", x"DD", x"77", -- 0x06B8,
      x"F6", x"DD", x"7E", x"F5", x"DD", x"77", x"F7", x"DD", -- 0x06C0,
      x"73", x"F8", x"DD", x"72", x"F9", x"AF", x"DD", x"77", -- 0x06C8,
      x"FF", x"DD", x"7E", x"F1", x"B7", x"28", x"10", x"0E", -- 0x06D0,
      x"03", x"DD", x"6E", x"F8", x"DD", x"66", x"F9", x"7E", -- 0x06D8,
      x"C6", x"E3", x"DD", x"77", x"FA", x"18", x"1F", x"DD", -- 0x06E0,
      x"6E", x"F2", x"DD", x"66", x"F3", x"7E", x"C6", x"E3", -- 0x06E8,
      x"4F", x"DD", x"6E", x"F6", x"DD", x"66", x"F7", x"7E", -- 0x06F0,
      x"B7", x"20", x"06", x"DD", x"36", x"FA", x"03", x"18", -- 0x06F8,
      x"05", x"C6", x"E3", x"DD", x"77", x"FA", x"26", x"00", -- 0x0700,
      x"69", x"29", x"29", x"29", x"DD", x"4E", x"FF", x"06", -- 0x0708,
      x"00", x"09", x"DD", x"75", x"FB", x"DD", x"74", x"FC", -- 0x0710,
      x"DD", x"6E", x"FA", x"26", x"00", x"29", x"29", x"29", -- 0x0718,
      x"09", x"4D", x"44", x"DD", x"7E", x"FB", x"C6", x"AF", -- 0x0720,
      x"6F", x"DD", x"7E", x"FC", x"CE", x"14", x"67", x"7E", -- 0x0728,
      x"87", x"87", x"87", x"87", x"DD", x"77", x"FC", x"21", -- 0x0730,
      x"AF", x"14", x"09", x"7E", x"07", x"07", x"07", x"07", -- 0x0738,
      x"E6", x"0F", x"DD", x"4E", x"FC", x"B1", x"D3", x"BE", -- 0x0740,
      x"DD", x"34", x"FF", x"DD", x"7E", x"FF", x"D6", x"08", -- 0x0748,
      x"DA", x"D1", x"06", x"DD", x"7E", x"FD", x"C6", x"10", -- 0x0750,
      x"DD", x"77", x"FD", x"30", x"03", x"DD", x"34", x"FE", -- 0x0758,
      x"DD", x"7E", x"F1", x"B7", x"28", x"07", x"AF", x"DD", -- 0x0760,
      x"77", x"F1", x"C3", x"9A", x"06", x"DD", x"5E", x"F4", -- 0x0768,
      x"DD", x"56", x"F5", x"C3", x"9A", x"06", x"DD", x"F9", -- 0x0770,
      x"DD", x"E1", x"C9", x"3E", x"8F", x"D3", x"BF", x"3E", -- 0x0778,
      x"AF", x"D3", x"BF", x"3E", x"00", x"D3", x"BE", x"3E", -- 0x0780,
      x"00", x"D3", x"BE", x"21", x"0A", x"00", x"E5", x"3E", -- 0x0788,
      x"F0", x"F5", x"33", x"21", x"03", x"10", x"E5", x"CD", -- 0x0790,
      x"46", x"37", x"F1", x"33", x"21", x"80", x"00", x"E3", -- 0x0798,
      x"21", x"4A", x"13", x"E5", x"21", x"40", x"02", x"E5", -- 0x07A0,
      x"CD", x"0A", x"29", x"F1", x"F1", x"F1", x"0E", x"01", -- 0x07A8,
      x"3E", x"8F", x"D3", x"BF", x"3E", x"AF", x"D3", x"BF", -- 0x07B0,
      x"79", x"D3", x"BE", x"79", x"87", x"87", x"87", x"87", -- 0x07B8,
      x"B1", x"D3", x"BE", x"C5", x"3E", x"03", x"F5", x"33", -- 0x07C0,
      x"CD", x"7A", x"02", x"33", x"C1", x"0C", x"79", x"D6", -- 0x07C8,
      x"10", x"38", x"DD", x"C9", x"CD", x"13", x"3F", x"F5", -- 0x07D0,
      x"21", x"13", x"00", x"E5", x"3E", x"60", x"F5", x"33", -- 0x07D8,
      x"21", x"0D", x"10", x"E5", x"CD", x"46", x"37", x"F1", -- 0x07E0,
      x"F1", x"33", x"01", x"3D", x"12", x"DD", x"36", x"FF", -- 0x07E8,
      x"10", x"C5", x"3E", x"02", x"F5", x"33", x"CD", x"7A", -- 0x07F0,
      x"02", x"33", x"C1", x"DD", x"6E", x"FF", x"26", x"00", -- 0x07F8,
      x"2B", x"29", x"29", x"29", x"29", x"29", x"EB", x"0A", -- 0x0800,
      x"03", x"6F", x"26", x"00", x"19", x"EB", x"0A", x"DD", -- 0x0808,
      x"77", x"FE", x"03", x"DD", x"6E", x"FE", x"26", x"00", -- 0x0810,
      x"C5", x"E5", x"C5", x"D5", x"CD", x"0A", x"29", x"F1", -- 0x0818,
      x"F1", x"F1", x"C1", x"79", x"DD", x"86", x"FE", x"4F", -- 0x0820,
      x"30", x"01", x"04", x"DD", x"35", x"FF", x"DD", x"7E", -- 0x0828,
      x"FF", x"B7", x"20", x"BD", x"F1", x"DD", x"E1", x"C9", -- 0x0830,
      x"CD", x"13", x"3F", x"F5", x"DD", x"6E", x"04", x"26", -- 0x0838,
      x"00", x"29", x"29", x"29", x"DD", x"75", x"FE", x"7C", -- 0x0840,
      x"C6", x"18", x"DD", x"77", x"FF", x"DD", x"4E", x"05", -- 0x0848,
      x"DD", x"46", x"06", x"59", x"50", x"1A", x"B7", x"28", -- 0x0850,
      x"1C", x"13", x"7B", x"4F", x"DD", x"96", x"05", x"6F", -- 0x0858,
      x"7A", x"DD", x"9E", x"06", x"67", x"3E", x"1F", x"BD", -- 0x0860,
      x"3E", x"00", x"9C", x"E2", x"70", x"08", x"EE", x"80", -- 0x0868,
      x"F2", x"55", x"08", x"AF", x"12", x"79", x"DD", x"4E", -- 0x0870,
      x"05", x"91", x"4F", x"41", x"2E", x"00", x"58", x"55", -- 0x0878,
      x"CB", x"7D", x"28", x"03", x"58", x"55", x"13", x"CB", -- 0x0880,
      x"2A", x"CB", x"1B", x"21", x"10", x"00", x"BF", x"ED", -- 0x0888,
      x"52", x"29", x"29", x"29", x"29", x"D1", x"D5", x"19", -- 0x0890,
      x"CB", x"41", x"28", x"15", x"01", x"F0", x"FF", x"09", -- 0x0898,
      x"4D", x"44", x"DD", x"6E", x"05", x"DD", x"66", x"06", -- 0x08A0,
      x"E5", x"C5", x"CD", x"7C", x"06", x"F1", x"F1", x"18", -- 0x08A8,
      x"0D", x"DD", x"4E", x"05", x"DD", x"46", x"06", x"C5", -- 0x08B0,
      x"E5", x"CD", x"35", x"06", x"F1", x"F1", x"F1", x"DD", -- 0x08B8,
      x"E1", x"C9", x"CD", x"13", x"3F", x"3B", x"3A", x"47", -- 0x08C0,
      x"73", x"E6", x"04", x"32", x"47", x"73", x"CD", x"1D", -- 0x08C8,
      x"14", x"3A", x"44", x"73", x"B7", x"28", x"13", x"01", -- 0x08D0,
      x"00", x"60", x"69", x"60", x"36", x"FF", x"23", x"36", -- 0x08D8,
      x"00", x"03", x"03", x"78", x"D6", x"64", x"38", x"F2", -- 0x08E0,
      x"18", x"10", x"01", x"00", x"60", x"59", x"50", x"AF", -- 0x08E8,
      x"12", x"13", x"12", x"03", x"03", x"78", x"D6", x"64", -- 0x08F0,
      x"38", x"F3", x"3A", x"00", x"80", x"D6", x"AA", x"C2", -- 0x08F8,
      x"EF", x"09", x"21", x"C8", x"63", x"36", x"33", x"3E", -- 0x0900,
      x"FF", x"D3", x"C0", x"21", x"08", x"80", x"4E", x"23", -- 0x0908,
      x"46", x"03", x"03", x"CB", x"A0", x"59", x"78", x"57", -- 0x0910,
      x"B1", x"28", x"0E", x"21", x"0A", x"00", x"E5", x"2E", -- 0x0918,
      x"00", x"E5", x"D5", x"CD", x"D1", x"00", x"F1", x"F1", -- 0x0920,
      x"F1", x"21", x"14", x"00", x"E5", x"2E", x"00", x"E5", -- 0x0928,
      x"21", x"07", x"63", x"E5", x"CD", x"D1", x"00", x"F1", -- 0x0930,
      x"F1", x"F1", x"21", x"06", x"00", x"E5", x"2E", x"00", -- 0x0938,
      x"E5", x"21", x"EB", x"63", x"E5", x"CD", x"D1", x"00", -- 0x0940,
      x"F1", x"F1", x"F1", x"21", x"C6", x"63", x"36", x"00", -- 0x0948,
      x"2E", x"C7", x"36", x"00", x"21", x"00", x"40", x"E5", -- 0x0950,
      x"AF", x"F5", x"33", x"26", x"00", x"E5", x"CD", x"46", -- 0x0958,
      x"37", x"F1", x"F1", x"33", x"DB", x"BF", x"DD", x"77", -- 0x0960,
      x"FF", x"3E", x"00", x"D3", x"BF", x"3E", x"80", x"D3", -- 0x0968,
      x"BF", x"21", x"C3", x"63", x"36", x"00", x"3E", x"80", -- 0x0970,
      x"D3", x"BF", x"3E", x"81", x"D3", x"BF", x"2E", x"C4", -- 0x0978,
      x"36", x"80", x"3E", x"06", x"D3", x"BF", x"3E", x"82", -- 0x0980,
      x"D3", x"BF", x"3E", x"80", x"D3", x"BF", x"3E", x"83", -- 0x0988,
      x"D3", x"BF", x"3E", x"00", x"D3", x"BF", x"3E", x"84", -- 0x0990,
      x"D3", x"BF", x"3E", x"36", x"D3", x"BF", x"3E", x"85", -- 0x0998,
      x"D3", x"BF", x"3E", x"07", x"D3", x"BF", x"3E", x"86", -- 0x09A0,
      x"D3", x"BF", x"21", x"0A", x"00", x"E5", x"21", x"B3", -- 0x09A8,
      x"01", x"E5", x"21", x"F2", x"63", x"E5", x"CD", x"AE", -- 0x09B0,
      x"00", x"F1", x"F1", x"21", x"00", x"03", x"E3", x"21", -- 0x09B8,
      x"AF", x"14", x"E5", x"21", x"E8", x"00", x"E5", x"CD", -- 0x09C0,
      x"0A", x"29", x"F1", x"F1", x"21", x"08", x"00", x"E3", -- 0x09C8,
      x"21", x"C7", x"14", x"E5", x"21", x"00", x"00", x"E5", -- 0x09D0,
      x"CD", x"0A", x"29", x"F1", x"F1", x"21", x"0F", x"00", -- 0x09D8,
      x"E3", x"21", x"A4", x"01", x"E5", x"21", x"03", x"20", -- 0x09E0,
      x"E5", x"CD", x"0A", x"29", x"F1", x"F1", x"F1", x"21", -- 0x09E8,
      x"09", x"00", x"E5", x"21", x"BD", x"01", x"E5", x"21", -- 0x09F0,
      x"00", x"60", x"E5", x"CD", x"AE", x"00", x"F1", x"F1", -- 0x09F8,
      x"F1", x"CD", x"00", x"60", x"33", x"DD", x"E1", x"C9", -- 0x0A00,
      x"3E", x"30", x"D3", x"55", x"C3", x"C2", x"08", x"CD", -- 0x0A08,
      x"13", x"3F", x"F5", x"F5", x"CD", x"B1", x"05", x"3A", -- 0x0A10,
      x"39", x"72", x"D6", x"12", x"20", x"03", x"CD", x"08", -- 0x0A18,
      x"0A", x"21", x"41", x"00", x"E5", x"2E", x"00", x"E5", -- 0x0A20,
      x"21", x"00", x"64", x"E5", x"CD", x"D1", x"00", x"F1", -- 0x0A28,
      x"F1", x"F1", x"1E", x"20", x"01", x"24", x"80", x"0A", -- 0x0A30,
      x"D6", x"2F", x"28", x"06", x"1D", x"28", x"03", x"03", -- 0x0A38,
      x"18", x"F5", x"7B", x"B7", x"20", x"05", x"C5", x"CD", -- 0x0A40,
      x"08", x"0A", x"C1", x"03", x"1E", x"20", x"0A", x"D6", -- 0x0A48,
      x"20", x"20", x"06", x"1D", x"28", x"03", x"03", x"18", -- 0x0A50,
      x"F5", x"11", x"38", x"0C", x"1A", x"DD", x"77", x"FE", -- 0x0A58,
      x"B7", x"28", x"10", x"0A", x"DD", x"77", x"FF", x"DD", -- 0x0A60,
      x"7E", x"FE", x"DD", x"96", x"FF", x"20", x"04", x"03", -- 0x0A68,
      x"13", x"18", x"E9", x"1E", x"20", x"0A", x"D6", x"20", -- 0x0A70,
      x"20", x"06", x"1D", x"28", x"03", x"03", x"18", x"F5", -- 0x0A78,
      x"DD", x"36", x"FD", x"20", x"11", x"00", x"64", x"0A", -- 0x0A80,
      x"6F", x"7B", x"C6", x"01", x"DD", x"77", x"FE", x"7A", -- 0x0A88,
      x"CE", x"00", x"DD", x"77", x"FF", x"7D", x"D6", x"2F", -- 0x0A90,
      x"28", x"14", x"DD", x"35", x"FD", x"DD", x"7E", x"FD", -- 0x0A98,
      x"B7", x"28", x"0B", x"7D", x"03", x"12", x"DD", x"5E", -- 0x0AA0,
      x"FE", x"DD", x"56", x"FF", x"18", x"D9", x"33", x"33", -- 0x0AA8,
      x"C5", x"3E", x"20", x"12", x"0E", x"20", x"11", x"24", -- 0x0AB0,
      x"80", x"1A", x"D6", x"20", x"20", x"06", x"0D", x"28", -- 0x0AB8,
      x"03", x"13", x"18", x"F5", x"DD", x"7E", x"FE", x"0E", -- 0x0AC0,
      x"00", x"91", x"4F", x"3E", x"39", x"91", x"4F", x"1A", -- 0x0AC8,
      x"47", x"D6", x"2F", x"28", x"15", x"0D", x"28", x"12", -- 0x0AD0,
      x"13", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"70", -- 0x0AD8,
      x"DD", x"34", x"FE", x"20", x"EA", x"DD", x"34", x"FF", -- 0x0AE0,
      x"18", x"E5", x"D1", x"C1", x"C5", x"D5", x"DD", x"36", -- 0x0AE8,
      x"FF", x"20", x"D1", x"D5", x"1A", x"13", x"D6", x"2F", -- 0x0AF0,
      x"3E", x"01", x"28", x"01", x"AF", x"6F", x"CB", x"45", -- 0x0AF8,
      x"20", x"09", x"DD", x"35", x"FF", x"DD", x"7E", x"FF", -- 0x0B00,
      x"B7", x"20", x"E9", x"7D", x"B7", x"28", x"19", x"3E", -- 0x0B08,
      x"20", x"02", x"03", x"3E", x"1D", x"02", x"03", x"1A", -- 0x0B10,
      x"13", x"02", x"03", x"1A", x"13", x"02", x"03", x"1A", -- 0x0B18,
      x"13", x"02", x"03", x"1A", x"02", x"03", x"AF", x"02", -- 0x0B20,
      x"0B", x"59", x"50", x"7B", x"D6", x"00", x"7A", x"DE", -- 0x0B28,
      x"64", x"38", x"09", x"0A", x"B7", x"20", x"F1", x"3E", -- 0x0B30,
      x"20", x"02", x"18", x"EC", x"21", x"40", x"64", x"36", -- 0x0B38,
      x"00", x"3A", x"00", x"64", x"D6", x"20", x"20", x"14", -- 0x0B40,
      x"21", x"40", x"00", x"E5", x"21", x"01", x"64", x"E5", -- 0x0B48,
      x"21", x"00", x"64", x"E5", x"CD", x"0B", x"01", x"F1", -- 0x0B50,
      x"F1", x"F1", x"18", x"E5", x"01", x"00", x"64", x"0A", -- 0x0B58,
      x"B7", x"28", x"39", x"59", x"50", x"13", x"D6", x"20", -- 0x0B60,
      x"20", x"2E", x"1A", x"D6", x"20", x"20", x"29", x"79", -- 0x0B68,
      x"D6", x"00", x"6F", x"78", x"DE", x"64", x"67", x"3E", -- 0x0B70,
      x"40", x"95", x"6F", x"3E", x"00", x"9C", x"67", x"DD", -- 0x0B78,
      x"71", x"FE", x"DD", x"70", x"FF", x"C5", x"E5", x"D5", -- 0x0B80,
      x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"E5", x"CD", -- 0x0B88,
      x"0B", x"01", x"F1", x"F1", x"F1", x"C1", x"18", x"C7", -- 0x0B90,
      x"4B", x"42", x"18", x"C3", x"11", x"40", x"64", x"4B", -- 0x0B98,
      x"42", x"79", x"D6", x"00", x"78", x"DE", x"64", x"38", -- 0x0BA0,
      x"07", x"1A", x"B7", x"20", x"03", x"1B", x"18", x"EF", -- 0x0BA8,
      x"7B", x"D6", x"00", x"4F", x"7A", x"DE", x"64", x"47", -- 0x0BB0,
      x"3E", x"1F", x"B9", x"3E", x"00", x"98", x"E2", x"C3", -- 0x0BB8,
      x"0B", x"EE", x"80", x"F2", x"04", x"0C", x"11", x"1E", -- 0x0BC0,
      x"64", x"4B", x"42", x"1A", x"D6", x"20", x"3E", x"01", -- 0x0BC8,
      x"28", x"01", x"AF", x"6F", x"3E", x"00", x"91", x"3E", -- 0x0BD0,
      x"64", x"98", x"30", x"07", x"CB", x"45", x"20", x"03", -- 0x0BD8,
      x"1B", x"18", x"E6", x"7D", x"B7", x"28", x"2A", x"AF", -- 0x0BE0,
      x"12", x"D5", x"21", x"00", x"64", x"E5", x"AF", x"F5", -- 0x0BE8,
      x"33", x"CD", x"38", x"08", x"F1", x"33", x"D1", x"13", -- 0x0BF0,
      x"D5", x"3E", x"01", x"F5", x"33", x"CD", x"38", x"08", -- 0x0BF8,
      x"F1", x"33", x"18", x"0D", x"21", x"00", x"64", x"E5", -- 0x0C00,
      x"3E", x"01", x"F5", x"33", x"CD", x"38", x"08", x"F1", -- 0x0C08,
      x"33", x"0E", x"FF", x"79", x"0D", x"B7", x"28", x"18", -- 0x0C10,
      x"C5", x"CD", x"B1", x"05", x"C1", x"3A", x"39", x"72", -- 0x0C18,
      x"D6", x"12", x"28", x"0C", x"C5", x"3E", x"01", x"F5", -- 0x0C20,
      x"33", x"CD", x"7A", x"02", x"33", x"C1", x"18", x"E3", -- 0x0C28,
      x"CD", x"08", x"0A", x"DD", x"F9", x"DD", x"E1", x"C9", -- 0x0C30,
      x"50", x"52", x"45", x"53", x"45", x"4E", x"54", x"53", -- 0x0C38,
      x"00", x"3B", x"E5", x"21", x"43", x"73", x"CB", x"86", -- 0x0C40,
      x"E1", x"21", x"00", x"40", x"E5", x"AF", x"F5", x"33", -- 0x0C48,
      x"26", x"00", x"E5", x"CD", x"46", x"37", x"F1", x"F1", -- 0x0C50,
      x"33", x"0E", x"00", x"79", x"D3", x"50", x"3E", x"00", -- 0x0C58,
      x"D3", x"51", x"0C", x"79", x"D6", x"10", x"38", x"F3", -- 0x0C60,
      x"CD", x"FB", x"13", x"CD", x"CA", x"13", x"3E", x"20", -- 0x0C68,
      x"D3", x"BF", x"3E", x"9E", x"D3", x"BF", x"3E", x"02", -- 0x0C70,
      x"F5", x"33", x"CD", x"56", x"01", x"33", x"FD", x"21", -- 0x0C78,
      x"00", x"00", x"FD", x"39", x"FD", x"75", x"00", x"3E", -- 0x0C80,
      x"00", x"D3", x"BF", x"3E", x"07", x"F6", x"40", x"D3", -- 0x0C88,
      x"BF", x"0E", x"00", x"3E", x"AF", x"D3", x"BE", x"79", -- 0x0C90,
      x"87", x"87", x"87", x"87", x"D3", x"BE", x"79", x"87", -- 0x0C98,
      x"87", x"D3", x"BE", x"3E", x"0F", x"D3", x"BE", x"0C", -- 0x0CA0,
      x"79", x"D6", x"10", x"38", x"E6", x"3E", x"D0", x"D3", -- 0x0CA8,
      x"BE", x"21", x"00", x"03", x"E5", x"3E", x"18", x"F5", -- 0x0CB0,
      x"33", x"26", x"00", x"E5", x"CD", x"46", x"37", x"F1", -- 0x0CB8,
      x"33", x"21", x"20", x"00", x"E3", x"3E", x"F0", x"F5", -- 0x0CC0,
      x"33", x"21", x"00", x"10", x"E5", x"CD", x"46", x"37", -- 0x0CC8,
      x"F1", x"33", x"21", x"13", x"05", x"E3", x"21", x"2A", -- 0x0CD0,
      x"0D", x"E5", x"21", x"00", x"08", x"E5", x"CD", x"C6", -- 0x0CD8,
      x"01", x"F1", x"F1", x"F1", x"21", x"00", x"00", x"39", -- 0x0CE0,
      x"7E", x"D3", x"BF", x"3E", x"81", x"D3", x"BF", x"3E", -- 0x0CE8,
      x"02", x"F5", x"33", x"CD", x"7A", x"02", x"33", x"3A", -- 0x0CF0,
      x"00", x"80", x"D6", x"55", x"20", x"0D", x"3A", x"01", -- 0x0CF8,
      x"80", x"D6", x"AA", x"20", x"06", x"CD", x"B1", x"05", -- 0x0D00,
      x"CD", x"08", x"0A", x"CD", x"7B", x"07", x"CD", x"D4", -- 0x0D08,
      x"07", x"21", x"00", x"80", x"7E", x"D6", x"AA", x"20", -- 0x0D10,
      x"0B", x"21", x"01", x"80", x"7E", x"D6", x"55", x"20", -- 0x0D18,
      x"03", x"CD", x"0F", x"0A", x"33", x"C3", x"5D", x"24", -- 0x0D20,
      x"33", x"C9", x"C0", x"7E", x"85", x"18", x"00", x"85", -- 0x0D28,
      x"C6", x"C2", x"7C", x"00", x"FC", x"82", x"C6", x"CB", -- 0x0D30,
      x"FC", x"CC", x"C6", x"00", x"7C", x"C6", x"C0", x"7C", -- 0x0D38,
      x"06", x"C6", x"7C", x"00", x"86", x"18", x"08", x"82", -- 0x0D40,
      x"C6", x"C5", x"D6", x"FE", x"EE", x"C6", x"00", x"7C", -- 0x0D48,
      x"82", x"C6", x"CA", x"FE", x"C6", x"C6", x"00", x"7C", -- 0x0D50,
      x"C6", x"C0", x"7C", x"06", x"C6", x"7C", x"08", x"82", -- 0x0D58,
      x"C6", x"C0", x"FE", x"82", x"C6", x"C9", x"00", x"FE", -- 0x0D60,
      x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"FC", -- 0x0D68,
      x"82", x"C6", x"CD", x"FC", x"CC", x"C6", x"00", x"FE", -- 0x0D70,
      x"C0", x"C0", x"FC", x"C0", x"C0", x"FE", x"00", x"07", -- 0x0D78,
      x"01", x"02", x"C4", x"11", x"0F", x"07", x"C0", x"E0", -- 0x0D80,
      x"83", x"F0", x"C5", x"E0", x"C0", x"FE", x"C0", x"C0", -- 0x0D88,
      x"FC", x"82", x"C0", x"C1", x"00", x"7C", x"84", x"C6", -- 0x0D90,
      x"C2", x"7C", x"00", x"FC", x"82", x"C6", x"C2", x"FC", -- 0x0D98,
      x"CC", x"C6", x"08", x"85", x"60", x"C1", x"7E", x"00", -- 0x0DA0,
      x"85", x"C6", x"CA", x"7C", x"00", x"C6", x"E6", x"F6", -- 0x0DA8,
      x"DE", x"CE", x"C6", x"C6", x"00", x"7C", x"82", x"C6", -- 0x0DB0,
      x"C2", x"FE", x"C6", x"C6", x"08", x"46", x"C0", x"80", -- 0x0DB8,
      x"46", x"C1", x"00", x"FE", x"45", x"C5", x"7F", x"07", -- 0x0DC0,
      x"07", x"87", x"C7", x"C7", x"82", x"E7", x"87", x"FE", -- 0x0DC8,
      x"88", x"01", x"C2", x"87", x"87", x"8F", x"83", x"9F", -- 0x0DD0,
      x"4E", x"C2", x"F0", x"F8", x"FE", x"45", x"82", x"0F", -- 0x0DD8,
      x"C1", x"8F", x"8F", x"82", x"CF", x"46", x"86", x"FC", -- 0x0DE0,
      x"C1", x"F8", x"00", x"46", x"C4", x"0F", x"81", x"E1", -- 0x0DE8,
      x"F1", x"F1", x"83", x"F9", x"C4", x"8F", x"87", x"83", -- 0x0DF0,
      x"81", x"81", x"82", x"80", x"C0", x"FE", x"44", x"CF", -- 0x0DF8,
      x"7F", x"3F", x"00", x"00", x"80", x"80", x"C0", x"E0", -- 0x0E00,
      x"F0", x"F9", x"07", x"0F", x"1F", x"3F", x"7F", x"7F", -- 0x0E08,
      x"42", x"C6", x"FE", x"FC", x"F8", x"F0", x"E0", x"E0", -- 0x0E10,
      x"C0", x"42", x"84", x"80", x"42", x"04", x"C2", x"FF", -- 0x0E18,
      x"FF", x"FC", x"04", x"C0", x"87", x"86", x"07", x"42", -- 0x0E20,
      x"84", x"FE", x"42", x"84", x"01", x"87", x"9F", x"85", -- 0x0E28,
      x"F0", x"41", x"05", x"41", x"85", x"7F", x"41", x"87", -- 0x0E30,
      x"CF", x"41", x"83", x"FC", x"43", x"03", x"C3", x"FF", -- 0x0E38,
      x"FF", x"F0", x"F0", x"03", x"C1", x"F8", x"FC", x"87", -- 0x0E40,
      x"80", x"87", x"0F", x"87", x"F9", x"86", x"80", x"C6", -- 0x0E48,
      x"81", x"07", x"0F", x"1F", x"1F", x"3F", x"7F", x"45", -- 0x0E50,
      x"C3", x"F9", x"F1", x"F0", x"E0", x"02", x"C4", x"80", -- 0x0E58,
      x"C0", x"E0", x"E0", x"F0", x"83", x"80", x"43", x"03", -- 0x0E60,
      x"43", x"83", x"7F", x"43", x"85", x"E7", x"C1", x"C7", -- 0x0E68,
      x"C7", x"83", x"FE", x"43", x"83", x"01", x"43", x"87", -- 0x0E70,
      x"F0", x"87", x"7F", x"82", x"FC", x"44", x"02", x"44", -- 0x0E78,
      x"02", x"C0", x"E0", x"83", x"F0", x"CB", x"1F", x"0F", -- 0x0E80,
      x"07", x"07", x"03", x"01", x"01", x"03", x"FF", x"FF", -- 0x0E88,
      x"FE", x"FC", x"82", x"F8", x"C1", x"FC", x"80", x"06", -- 0x0E90,
      x"44", x"02", x"84", x"80", x"02", x"84", x"07", x"02", -- 0x0E98,
      x"83", x"FE", x"C0", x"FC", x"02", x"84", x"01", x"02", -- 0x0EA0,
      x"C4", x"9F", x"8F", x"8F", x"87", x"01", x"02", x"42", -- 0x0EA8,
      x"C1", x"FE", x"FC", x"02", x"C3", x"87", x"87", x"03", -- 0x0EB0,
      x"01", x"03", x"43", x"C0", x"7F", x"02", x"83", x"FC", -- 0x0EB8,
      x"C0", x"F8", x"02", x"84", x"0F", x"02", x"84", x"F9", -- 0x0EC0,
      x"02", x"C4", x"81", x"83", x"87", x"8F", x"8F", x"02", -- 0x0EC8,
      x"43", x"C0", x"FE", x"02", x"C2", x"C0", x"80", x"80", -- 0x0ED0,
      x"04", x"C4", x"3F", x"3F", x"1F", x"0F", x"07", x"02", -- 0x0ED8,
      x"C4", x"F8", x"FC", x"FE", x"FE", x"FF", x"02", x"77", -- 0x0EE0,
      x"07", x"C2", x"3F", x"7F", x"7F", x"84", x"3F", x"C1", -- 0x0EE8,
      x"FE", x"FE", x"45", x"03", x"C3", x"80", x"F0", x"FC", -- 0x0EF0,
      x"FC", x"04", x"C2", x"01", x"01", x"07", x"4A", x"84", -- 0x0EF8,
      x"FE", x"C0", x"80", x"06", x"C0", x"7F", x"86", x"3F", -- 0x0F00,
      x"C7", x"83", x"81", x"C1", x"C1", x"A0", x"A0", x"80", -- 0x0F08,
      x"C0", x"84", x"F8", x"C2", x"FC", x"7C", x"7C", x"05", -- 0x0F10,
      x"C1", x"01", x"01", x"02", x"C5", x"01", x"03", x"8F", -- 0x0F18,
      x"FF", x"FF", x"7F", x"46", x"C2", x"F0", x"F8", x"FC", -- 0x0F20,
      x"44", x"C2", x"00", x"00", x"7E", x"44", x"04", x"C2", -- 0x0F28,
      x"80", x"C0", x"C0", x"03", x"C5", x"01", x"03", x"0F", -- 0x0F30,
      x"1F", x"3F", x"7F", x"42", x"CA", x"FE", x"FC", x"F8", -- 0x0F38,
      x"F0", x"E0", x"C0", x"C1", x"80", x"00", x"01", x"01", -- 0x0F40,
      x"02", x"C4", x"80", x"F0", x"F0", x"E0", x"E0", x"83", -- 0x0F48,
      x"0F", x"83", x"07", x"D1", x"F0", x"F8", x"F8", x"FC", -- 0x0F50,
      x"FE", x"F9", x"E1", x"E0", x"F0", x"78", x"28", x"14", -- 0x0F58,
      x"08", x"04", x"80", x"C0", x"03", x"01", x"05", x"42", -- 0x0F60,
      x"C5", x"1F", x"0F", x"03", x"01", x"00", x"8F", x"4D", -- 0x0F68,
      x"CB", x"FE", x"FE", x"F8", x"F0", x"E0", x"C0", x"80", -- 0x0F70,
      x"00", x"00", x"03", x"07", x"07", x"03", x"CB", x"01", -- 0x0F78,
      x"F0", x"C1", x"03", x"07", x"0F", x"3F", x"FF", x"FF", -- 0x0F80,
      x"F8", x"F9", x"F9", x"49", x"C7", x"FE", x"FE", x"FC", -- 0x0F88,
      x"FE", x"FE", x"FC", x"98", x"10", x"02", x"C7", x"33", -- 0x0F90,
      x"40", x"80", x"00", x"00", x"01", x"03", x"07", x"83", -- 0x0F98,
      x"7F", x"43", x"C1", x"F0", x"FC", x"45", x"C2", x"1F", -- 0x0FA0,
      x"1F", x"0F", x"82", x"1F", x"C5", x"01", x"00", x"FE", -- 0x0FA8,
      x"FF", x"FE", x"FE", x"43", x"C8", x"60", x"30", x"98", -- 0x0FB0,
      x"4C", x"22", x"80", x"C0", x"80", x"07", x"06", x"C0", -- 0x0FB8,
      x"10", x"06", x"C1", x"1F", x"1C", x"05", x"C0", x"E0", -- 0x0FC0,
      x"0B", x"C7", x"01", x"07", x"1F", x"05", x"03", x"07", -- 0x0FC8,
      x"1F", x"7F", x"42", x"C1", x"C0", x"C0", x"82", x"80", -- 0x0FD0,
      x"02", x"86", x"01", x"C8", x"00", x"FE", x"FC", x"FE", -- 0x0FD8,
      x"FC", x"FE", x"FF", x"FF", x"1F", x"02", x"C4", x"08", -- 0x0FE0,
      x"01", x"80", x"C0", x"F8", x"04", x"C0", x"20", x"06", -- 0x0FE8,
      x"CA", x"07", x"00", x"00", x"1E", x"78", x"07", x"1F", -- 0x0FF0,
      x"FF", x"8F", x"1F", x"E7", x"44", x"C6", x"FE", x"FC", -- 0x0FF8,
      x"F8", x"80", x"C0", x"80", x"80", x"03", x"83", x"07", -- 0x1000,
      x"C4", x"0F", x"0F", x"06", x"00", x"FC", x"44", x"C3", -- 0x1008,
      x"7F", x"7F", x"00", x"00", x"45", x"02", x"C4", x"F8", -- 0x1010,
      x"F8", x"F0", x"F8", x"F8", x"02", x"C4", x"04", x"06", -- 0x1018,
      x"07", x"07", x"03", x"04", x"C6", x"81", x"F1", x"FF", -- 0x1020,
      x"00", x"00", x"F0", x"FE", x"43", x"C3", x"0F", x"0F", -- 0x1028,
      x"7F", x"3F", x"48", x"C2", x"F1", x"C0", x"80", x"43", -- 0x1030,
      x"CC", x"F1", x"E0", x"00", x"00", x"FE", x"FE", x"FC", -- 0x1038,
      x"F8", x"F8", x"F0", x"00", x"00", x"3C", x"06", x"82", -- 0x1040,
      x"07", x"84", x"03", x"87", x"F0", x"03", x"C5", x"70", -- 0x1048,
      x"70", x"78", x"78", x"00", x"01", x"05", x"CA", x"C0", -- 0x1050,
      x"C0", x"D0", x"D0", x"D3", x"F3", x"FB", x"7B", x"FF", -- 0x1058,
      x"7F", x"7F", x"44", x"C0", x"C0", x"82", x"80", x"83", -- 0x1060,
      x"C0", x"C0", x"01", x"06", x"C7", x"FF", x"CF", x"0F", -- 0x1068,
      x"07", x"07", x"03", x"01", x"00", x"42", x"C7", x"FE", -- 0x1070,
      x"FC", x"F8", x"E0", x"00", x"FF", x"8F", x"07", x"04", -- 0x1078,
      x"C4", x"FF", x"FF", x"3F", x"1F", x"0F", x"03", x"82", -- 0x1080,
      x"80", x"08", x"C2", x"0F", x"0F", x"1F", x"03", x"C3", -- 0x1088,
      x"06", x"1E", x"FE", x"FE", x"02", x"C4", x"18", x"3E", -- 0x1090,
      x"7F", x"7F", x"FF", x"02", x"C1", x"04", x"0E", x"42", -- 0x1098,
      x"05", x"C3", x"C0", x"C0", x"3F", x"3F", x"84", x"7F", -- 0x10A0,
      x"C4", x"3F", x"FF", x"FF", x"CF", x"8F", x"82", x"C7", -- 0x10A8,
      x"C0", x"C3", x"84", x"FC", x"CA", x"FE", x"FE", x"FF", -- 0x10B0,
      x"00", x"00", x"08", x"0C", x"1C", x"3C", x"7E", x"7F", -- 0x10B8,
      x"06", x"C0", x"E0", x"82", x"3F", x"82", x"1F", x"C1", -- 0x10C0,
      x"3F", x"3F", x"45", x"C3", x"FC", x"F0", x"FE", x"FE", -- 0x10C8,
      x"83", x"FC", x"C2", x"7E", x"7E", x"0F", x"86", x"1F", -- 0x10D0,
      x"45", x"D5", x"F1", x"F0", x"C0", x"E0", x"E0", x"D0", -- 0x10D8,
      x"C0", x"E0", x"E0", x"F0", x"3E", x"3F", x"1F", x"1F", -- 0x10E0,
      x"0F", x"0F", x"07", x"07", x"00", x"00", x"FC", x"FC", -- 0x10E8,
      x"82", x"FE", x"40", x"05", x"C0", x"01", x"84", x"03", -- 0x10F0,
      x"C2", x"07", x"07", x"0F", x"44", x"C7", x"FC", x"F0", -- 0x10F8,
      x"C0", x"00", x"FF", x"FF", x"FE", x"B8", x"02", x"C8", -- 0x1100,
      x"01", x"FF", x"87", x"03", x"0F", x"1F", x"7F", x"FF", -- 0x1108,
      x"FD", x"82", x"E0", x"83", x"F0", x"C0", x"F8", x"02", -- 0x1110,
      x"C7", x"01", x"1F", x"7F", x"FF", x"FF", x"1F", x"3F", -- 0x1118,
      x"7F", x"44", x"CF", x"F8", x"F0", x"F0", x"E0", x"C0", -- 0x1120,
      x"80", x"80", x"00", x"03", x"03", x"07", x"07", x"0F", -- 0x1128,
      x"0F", x"1F", x"3F", x"87", x"E0", x"C0", x"3F", x"44", -- 0x1130,
      x"EC", x"7F", x"3F", x"E0", x"F0", x"F8", x"FC", x"FE", -- 0x1138,
      x"FF", x"F9", x"FC", x"60", x"30", x"18", x"0C", x"06", -- 0x1140,
      x"00", x"80", x"C0", x"7F", x"3F", x"1F", x"0F", x"03", -- 0x1148,
      x"01", x"00", x"00", x"FC", x"F8", x"F9", x"FB", x"FF", -- 0x1150,
      x"3F", x"3F", x"0F", x"00", x"40", x"E0", x"F4", x"FC", -- 0x1158,
      x"FC", x"F8", x"F8", x"07", x"1F", x"7F", x"42", x"C1", -- 0x1160,
      x"DF", x"1F", x"45", x"C1", x"FE", x"F8", x"43", x"C7", -- 0x1168,
      x"FE", x"FC", x"F0", x"00", x"F8", x"E0", x"C0", x"80", -- 0x1170,
      x"03", x"CF", x"07", x"0F", x"1E", x"3C", x"78", x"01", -- 0x1178,
      x"01", x"02", x"FF", x"FF", x"7F", x"7F", x"FF", x"FF", -- 0x1180,
      x"BF", x"7F", x"44", x"C2", x"F3", x"F1", x"E1", x"82", -- 0x1188,
      x"80", x"82", x"C0", x"C4", x"80", x"80", x"FF", x"FF", -- 0x1190,
      x"03", x"84", x"01", x"82", x"80", x"C7", x"C0", x"E0", -- 0x1198,
      x"F8", x"FC", x"FE", x"00", x"01", x"01", x"04", x"C2", -- 0x11A0,
      x"FF", x"FF", x"81", x"02", x"CC", x"01", x"07", x"EF", -- 0x11A8,
      x"DF", x"3F", x"7F", x"7F", x"FF", x"BF", x"3F", x"FF", -- 0x11B0,
      x"FE", x"FE", x"44", x"06", x"C2", x"80", x"1F", x"1F", -- 0x11B8,
      x"82", x"0F", x"82", x"07", x"C3", x"FE", x"F7", x"F0", -- 0x11C0,
      x"F0", x"82", x"F8", x"C5", x"FC", x"30", x"86", x"00", -- 0x11C8,
      x"00", x"04", x"07", x"CC", x"06", x"00", x"07", x"1F", -- 0x11D0,
      x"38", x"03", x"3F", x"7F", x"3F", x"1F", x"FF", x"87", -- 0x11D8,
      x"1F", x"45", x"C1", x"F0", x"F0", x"82", x"E0", x"C2", -- 0x11E0,
      x"E3", x"FF", x"FF", x"83", x"3F", x"C3", x"3E", x"3E", -- 0x11E8,
      x"7E", x"7E", x"42", x"C5", x"7F", x"3F", x"1F", x"0F", -- 0x11F0,
      x"0F", x"E1", x"46", x"86", x"F8", x"C5", x"F0", x"03", -- 0x11F8,
      x"03", x"01", x"81", x"81", x"82", x"80", x"45", x"C5", -- 0x1200,
      x"E6", x"C6", x"FF", x"F1", x"C0", x"80", x"03", x"42", -- 0x1208,
      x"C1", x"FE", x"3C", x"02", x"82", x"03", x"C1", x"01", -- 0x1210,
      x"01", x"02", x"45", x"C5", x"3F", x"03", x"E0", x"E0", -- 0x1218,
      x"F8", x"F8", x"43", x"C4", x"78", x"F8", x"F9", x"FD", -- 0x1220,
      x"FD", x"42", x"C9", x"00", x"00", x"20", x"30", x"90", -- 0x1228,
      x"9C", x"FD", x"FF", x"7F", x"7F", x"46", x"82", x"FE", -- 0x1230,
      x"C3", x"FC", x"F8", x"F0", x"C0", x"0C", x"06", x"B2", -- 0x1238,
      x"B3", x"B4", x"B5", x"B6", x"B7", x"0B", x"07", x"F9", -- 0x1240,
      x"FA", x"FB", x"FC", x"FD", x"FE", x"FF", x"0A", x"09", -- 0x1248,
      x"AA", x"AB", x"6D", x"AC", x"AD", x"AE", x"AF", x"B0", -- 0x1250,
      x"B1", x"0A", x"0B", x"F1", x"F2", x"F3", x"F4", x"68", -- 0x1258,
      x"68", x"F5", x"6D", x"F6", x"F7", x"F8", x"09", x"0F", -- 0x1260,
      x"9F", x"A0", x"A1", x"A2", x"68", x"68", x"68", x"A3", -- 0x1268,
      x"A4", x"A5", x"A6", x"6D", x"A7", x"A8", x"A9", x"09", -- 0x1270,
      x"0F", x"EA", x"EB", x"68", x"68", x"68", x"68", x"68", -- 0x1278,
      x"68", x"68", x"68", x"ED", x"EE", x"EF", x"6D", x"F0", -- 0x1280,
      x"08", x"11", x"97", x"98", x"99", x"68", x"68", x"68", -- 0x1288,
      x"68", x"68", x"68", x"68", x"68", x"68", x"9B", x"9C", -- 0x1290,
      x"75", x"9D", x"9E", x"08", x"11", x"E3", x"E4", x"68", -- 0x1298,
      x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"68", -- 0x12A0,
      x"68", x"E5", x"E6", x"E7", x"E8", x"E9", x"07", x"12", -- 0x12A8,
      x"8D", x"8E", x"8F", x"68", x"68", x"68", x"90", x"91", -- 0x12B0,
      x"68", x"92", x"93", x"68", x"68", x"68", x"94", x"95", -- 0x12B8,
      x"6D", x"96", x"07", x"13", x"D5", x"D6", x"D7", x"68", -- 0x12C0,
      x"68", x"D8", x"D9", x"DA", x"68", x"DB", x"DC", x"DD", -- 0x12C8,
      x"DE", x"68", x"68", x"DF", x"E0", x"E1", x"E2", x"07", -- 0x12D0,
      x"12", x"7D", x"7E", x"7F", x"80", x"81", x"82", x"83", -- 0x12D8,
      x"84", x"68", x"85", x"86", x"87", x"88", x"89", x"68", -- 0x12E0,
      x"8A", x"8B", x"8C", x"07", x"12", x"C5", x"C6", x"C7", -- 0x12E8,
      x"C8", x"C9", x"CA", x"CB", x"6D", x"CC", x"CD", x"CE", -- 0x12F0,
      x"CF", x"D0", x"D1", x"D2", x"D3", x"6D", x"D4", x"08", -- 0x12F8,
      x"11", x"70", x"71", x"72", x"68", x"68", x"73", x"74", -- 0x1300,
      x"75", x"76", x"77", x"78", x"68", x"79", x"7A", x"7B", -- 0x1308,
      x"6A", x"7C", x"08", x"10", x"BD", x"BE", x"BF", x"68", -- 0x1310,
      x"68", x"68", x"68", x"C0", x"C1", x"68", x"68", x"68", -- 0x1318,
      x"68", x"C2", x"C3", x"C4", x"08", x"11", x"69", x"6A", -- 0x1320,
      x"6B", x"68", x"68", x"68", x"68", x"68", x"68", x"68", -- 0x1328,
      x"68", x"68", x"68", x"6C", x"6D", x"6E", x"6F", x"08", -- 0x1330,
      x"11", x"B8", x"B9", x"68", x"68", x"68", x"68", x"68", -- 0x1338,
      x"68", x"68", x"68", x"68", x"68", x"68", x"68", x"BA", -- 0x1340,
      x"BB", x"BC", x"18", x"20", x"19", x"1A", x"1B", x"1C", -- 0x1348,
      x"1D", x"18", x"1E", x"20", x"1F", x"21", x"1A", x"1A", -- 0x1350,
      x"22", x"23", x"24", x"1A", x"1A", x"25", x"20", x"19", -- 0x1358,
      x"1A", x"26", x"27", x"20", x"28", x"29", x"2A", x"2B", -- 0x1360,
      x"2C", x"18", x"18", x"20", x"42", x"43", x"44", x"45", -- 0x1368,
      x"46", x"43", x"47", x"20", x"33", x"48", x"18", x"18", -- 0x1370,
      x"49", x"37", x"4A", x"4B", x"4B", x"4C", x"20", x"3B", -- 0x1378,
      x"18", x"3C", x"3D", x"20", x"3B", x"4D", x"20", x"4E", -- 0x1380,
      x"4F", x"18", x"18", x"20", x"2D", x"2E", x"2F", x"30", -- 0x1388,
      x"31", x"2E", x"32", x"20", x"33", x"34", x"35", x"35", -- 0x1390,
      x"36", x"37", x"38", x"39", x"39", x"3A", x"20", x"3B", -- 0x1398,
      x"18", x"3C", x"3D", x"20", x"3E", x"3F", x"40", x"1B", -- 0x13A0,
      x"41", x"18", x"18", x"50", x"51", x"18", x"18", x"52", -- 0x13A8,
      x"53", x"18", x"54", x"50", x"55", x"50", x"50", x"50", -- 0x13B0,
      x"56", x"57", x"58", x"50", x"50", x"59", x"50", x"51", -- 0x13B8,
      x"18", x"5A", x"5B", x"50", x"5C", x"5D", x"5E", x"5F", -- 0x13C0,
      x"60", x"18", x"3E", x"1C", x"D3", x"BF", x"3E", x"B9", -- 0x13C8,
      x"D3", x"BF", x"3E", x"1C", x"D3", x"BF", x"3E", x"B9", -- 0x13D0,
      x"D3", x"BF", x"C9", x"00", x"00", x"00", x"00", x"C3", -- 0x13D8,
      x"02", x"D6", x"05", x"4F", x"05", x"6F", x"07", x"54", -- 0x13E0,
      x"0D", x"EF", x"04", x"54", x"0F", x"76", x"0F", x"C3", -- 0x13E8,
      x"0D", x"D6", x"0E", x"B2", x"02", x"5C", x"0C", x"CC", -- 0x13F0,
      x"0C", x"FF", x"0F", x"3E", x"80", x"D3", x"BF", x"3E", -- 0x13F8,
      x"B2", x"D3", x"BF", x"3E", x"00", x"D3", x"BF", x"3E", -- 0x1400,
      x"87", x"D3", x"BF", x"3E", x"80", x"D3", x"BF", x"3E", -- 0x1408,
      x"81", x"D3", x"BF", x"C9", x"3E", x"00", x"D3", x"BF", -- 0x1410,
      x"3E", x"B9", x"D3", x"BF", x"C9", x"CD", x"FB", x"13", -- 0x1418,
      x"CD", x"CA", x"13", x"3E", x"00", x"D3", x"BF", x"3E", -- 0x1420,
      x"B8", x"D3", x"BF", x"3E", x"00", x"D3", x"BF", x"3E", -- 0x1428,
      x"98", x"D3", x"BF", x"3E", x"10", x"F5", x"33", x"21", -- 0x1430,
      x"DB", x"13", x"E5", x"CD", x"7D", x"14", x"F1", x"33", -- 0x1438,
      x"3E", x"00", x"D3", x"BF", x"3E", x"8F", x"D3", x"BF", -- 0x1440,
      x"3A", x"45", x"73", x"B7", x"28", x"0A", x"3E", x"04", -- 0x1448,
      x"D3", x"BF", x"3E", x"9E", x"D3", x"BF", x"18", x"08", -- 0x1450,
      x"3E", x"20", x"D3", x"BF", x"3E", x"9E", x"D3", x"BF", -- 0x1458,
      x"FD", x"21", x"47", x"73", x"FD", x"7E", x"00", x"D3", -- 0x1460,
      x"BF", x"3E", x"B2", x"D3", x"BF", x"DB", x"BF", x"07", -- 0x1468,
      x"D2", x"14", x"14", x"00", x"00", x"00", x"00", x"00", -- 0x1470,
      x"18", x"F3", x"C3", x"14", x"14", x"CD", x"13", x"3F", -- 0x1478,
      x"3E", x"C0", x"D3", x"BF", x"3E", x"AF", x"D3", x"BF", -- 0x1480,
      x"DD", x"4E", x"04", x"DD", x"46", x"05", x"DD", x"5E", -- 0x1488,
      x"06", x"7B", x"1D", x"B7", x"28", x"0E", x"69", x"60", -- 0x1490,
      x"56", x"23", x"7E", x"D3", x"BE", x"0A", x"D3", x"BE", -- 0x1498,
      x"03", x"03", x"18", x"ED", x"3E", x"00", x"D3", x"BF", -- 0x14A0,
      x"3E", x"AF", x"D3", x"BF", x"DD", x"E1", x"C9", x"78", -- 0x14A8,
      x"84", x"B4", x"A4", x"B4", x"84", x"78", x"00", x"1F", -- 0x14B0,
      x"04", x"04", x"04", x"00", x"00", x"00", x"00", x"44", -- 0x14B8,
      x"6C", x"54", x"54", x"00", x"00", x"00", x"00", x"00", -- 0x14C0,
      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", -- 0x14C8,
      x"20", x"20", x"20", x"00", x"00", x"20", x"00", x"50", -- 0x14D0,
      x"50", x"50", x"00", x"00", x"00", x"00", x"00", x"50", -- 0x14D8,
      x"50", x"F8", x"50", x"F8", x"50", x"50", x"00", x"20", -- 0x14E0,
      x"78", x"A0", x"70", x"28", x"F0", x"20", x"00", x"C0", -- 0x14E8,
      x"C8", x"10", x"20", x"40", x"98", x"18", x"00", x"40", -- 0x14F0,
      x"A0", x"40", x"A8", x"90", x"98", x"60", x"00", x"10", -- 0x14F8,
      x"20", x"40", x"00", x"00", x"00", x"00", x"00", x"10", -- 0x1500,
      x"20", x"40", x"40", x"40", x"20", x"10", x"00", x"40", -- 0x1508,
      x"20", x"10", x"10", x"10", x"20", x"40", x"00", x"20", -- 0x1510,
      x"A8", x"70", x"20", x"70", x"A8", x"20", x"00", x"00", -- 0x1518,
      x"20", x"20", x"F8", x"20", x"20", x"00", x"00", x"00", -- 0x1520,
      x"00", x"00", x"00", x"00", x"20", x"20", x"40", x"00", -- 0x1528,
      x"00", x"00", x"78", x"00", x"00", x"00", x"00", x"00", -- 0x1530,
      x"00", x"00", x"00", x"00", x"60", x"60", x"00", x"00", -- 0x1538,
      x"00", x"08", x"10", x"20", x"40", x"80", x"00", x"70", -- 0x1540,
      x"88", x"98", x"A8", x"C8", x"88", x"70", x"00", x"20", -- 0x1548,
      x"60", x"20", x"20", x"20", x"20", x"70", x"00", x"70", -- 0x1550,
      x"88", x"08", x"10", x"60", x"80", x"F8", x"00", x"70", -- 0x1558,
      x"88", x"08", x"30", x"08", x"88", x"70", x"00", x"10", -- 0x1560,
      x"30", x"50", x"90", x"F8", x"10", x"10", x"00", x"F8", -- 0x1568,
      x"80", x"E0", x"10", x"08", x"10", x"E0", x"00", x"30", -- 0x1570,
      x"40", x"80", x"F0", x"88", x"88", x"70", x"00", x"F8", -- 0x1578,
      x"88", x"10", x"20", x"20", x"20", x"20", x"00", x"70", -- 0x1580,
      x"88", x"88", x"70", x"88", x"88", x"70", x"00", x"70", -- 0x1588,
      x"88", x"88", x"78", x"08", x"10", x"60", x"00", x"00", -- 0x1590,
      x"00", x"20", x"00", x"00", x"20", x"00", x"00", x"00", -- 0x1598,
      x"00", x"20", x"00", x"00", x"20", x"20", x"40", x"18", -- 0x15A0,
      x"30", x"60", x"C0", x"60", x"30", x"18", x"00", x"00", -- 0x15A8,
      x"00", x"F8", x"00", x"F8", x"00", x"00", x"00", x"C0", -- 0x15B0,
      x"60", x"30", x"18", x"30", x"60", x"C0", x"00", x"70", -- 0x15B8,
      x"88", x"08", x"10", x"20", x"00", x"20", x"00", x"70", -- 0x15C0,
      x"88", x"08", x"48", x"A8", x"A8", x"70", x"00", x"20", -- 0x15C8,
      x"50", x"88", x"88", x"F8", x"88", x"88", x"00", x"F0", -- 0x15D0,
      x"48", x"48", x"70", x"48", x"48", x"F0", x"00", x"30", -- 0x15D8,
      x"48", x"80", x"80", x"80", x"48", x"30", x"00", x"E0", -- 0x15E0,
      x"50", x"48", x"48", x"48", x"50", x"E0", x"00", x"F8", -- 0x15E8,
      x"80", x"80", x"F0", x"80", x"80", x"F8", x"00", x"F8", -- 0x15F0,
      x"80", x"80", x"F0", x"80", x"80", x"80", x"00", x"70", -- 0x15F8,
      x"88", x"80", x"B8", x"88", x"88", x"70", x"00", x"88", -- 0x1600,
      x"88", x"88", x"F8", x"88", x"88", x"88", x"00", x"70", -- 0x1608,
      x"20", x"20", x"20", x"20", x"20", x"70", x"00", x"38", -- 0x1610,
      x"10", x"10", x"10", x"90", x"90", x"60", x"00", x"88", -- 0x1618,
      x"90", x"A0", x"C0", x"A0", x"90", x"88", x"00", x"80", -- 0x1620,
      x"80", x"80", x"80", x"80", x"80", x"F8", x"00", x"88", -- 0x1628,
      x"D8", x"A8", x"A8", x"88", x"88", x"88", x"00", x"88", -- 0x1630,
      x"C8", x"C8", x"A8", x"98", x"98", x"88", x"00", x"70", -- 0x1638,
      x"88", x"88", x"88", x"88", x"88", x"70", x"00", x"F0", -- 0x1640,
      x"88", x"88", x"F0", x"80", x"80", x"80", x"00", x"70", -- 0x1648,
      x"88", x"88", x"88", x"A8", x"90", x"68", x"00", x"F0", -- 0x1650,
      x"88", x"88", x"F0", x"A0", x"90", x"88", x"00", x"70", -- 0x1658,
      x"88", x"80", x"70", x"08", x"88", x"70", x"00", x"F8", -- 0x1660,
      x"20", x"20", x"20", x"20", x"20", x"20", x"00", x"88", -- 0x1668,
      x"88", x"88", x"88", x"88", x"88", x"70", x"00", x"88", -- 0x1670,
      x"88", x"88", x"88", x"50", x"50", x"20", x"00", x"88", -- 0x1678,
      x"88", x"88", x"A8", x"A8", x"D8", x"88", x"00", x"88", -- 0x1680,
      x"88", x"50", x"20", x"50", x"88", x"88", x"00", x"88", -- 0x1688,
      x"88", x"88", x"70", x"20", x"20", x"20", x"00", x"F8", -- 0x1690,
      x"08", x"10", x"20", x"40", x"80", x"F8", x"00", x"70", -- 0x1698,
      x"40", x"40", x"40", x"40", x"40", x"70", x"00", x"00", -- 0x16A0,
      x"00", x"80", x"40", x"20", x"10", x"08", x"00", x"70", -- 0x16A8,
      x"10", x"10", x"10", x"10", x"10", x"70", x"00", x"20", -- 0x16B0,
      x"50", x"88", x"00", x"00", x"00", x"00", x"00", x"00", -- 0x16B8,
      x"00", x"00", x"00", x"00", x"00", x"F8", x"00", x"80", -- 0x16C0,
      x"40", x"20", x"00", x"00", x"00", x"00", x"00", x"00", -- 0x16C8,
      x"00", x"70", x"08", x"78", x"88", x"78", x"00", x"80", -- 0x16D0,
      x"80", x"B0", x"C8", x"88", x"C8", x"B0", x"00", x"00", -- 0x16D8,
      x"00", x"70", x"88", x"80", x"88", x"70", x"00", x"08", -- 0x16E0,
      x"08", x"68", x"98", x"88", x"98", x"68", x"00", x"00", -- 0x16E8,
      x"00", x"70", x"88", x"F8", x"80", x"70", x"00", x"10", -- 0x16F0,
      x"28", x"20", x"F8", x"20", x"20", x"20", x"00", x"00", -- 0x16F8,
      x"00", x"68", x"98", x"98", x"68", x"08", x"70", x"80", -- 0x1700,
      x"80", x"F0", x"88", x"88", x"88", x"88", x"00", x"20", -- 0x1708,
      x"00", x"60", x"20", x"20", x"20", x"70", x"00", x"10", -- 0x1710,
      x"00", x"30", x"10", x"10", x"10", x"90", x"60", x"40", -- 0x1718,
      x"40", x"48", x"50", x"60", x"50", x"48", x"00", x"60", -- 0x1720,
      x"20", x"20", x"20", x"20", x"20", x"70", x"00", x"00", -- 0x1728,
      x"00", x"D0", x"A8", x"A8", x"A8", x"A8", x"00", x"00", -- 0x1730,
      x"00", x"B0", x"C8", x"88", x"88", x"88", x"00", x"00", -- 0x1738,
      x"00", x"70", x"88", x"88", x"88", x"70", x"00", x"00", -- 0x1740,
      x"00", x"B0", x"C8", x"C8", x"B0", x"80", x"80", x"00", -- 0x1748,
      x"00", x"68", x"98", x"98", x"68", x"08", x"08", x"00", -- 0x1750,
      x"00", x"B0", x"C8", x"80", x"80", x"80", x"00", x"00", -- 0x1758,
      x"00", x"78", x"80", x"70", x"08", x"F0", x"00", x"40", -- 0x1760,
      x"40", x"F0", x"40", x"40", x"48", x"30", x"00", x"00", -- 0x1768,
      x"00", x"90", x"90", x"90", x"90", x"68", x"00", x"00", -- 0x1770,
      x"00", x"88", x"88", x"88", x"50", x"20", x"00", x"00", -- 0x1778,
      x"00", x"88", x"A8", x"A8", x"A8", x"50", x"00", x"00", -- 0x1780,
      x"00", x"88", x"50", x"20", x"50", x"88", x"00", x"00", -- 0x1788,
      x"00", x"88", x"88", x"98", x"68", x"08", x"70", x"00", -- 0x1790,
      x"00", x"F8", x"10", x"20", x"40", x"F8", x"00", x"FD", -- 0x1798,
      x"21", x"02", x"00", x"FD", x"39", x"FD", x"4E", x"00", -- 0x17A0,
      x"79", x"0D", x"B7", x"C8", x"E3", x"E3", x"E3", x"E3", -- 0x17A8,
      x"E3", x"E3", x"E3", x"E3", x"18", x"F2", x"43", x"4F", -- 0x17B0,
      x"4C", x"45", x"43", x"4F", x"00", x"07", x"00", x"00", -- 0x17B8,
      x"00", x"00", x"00", x"00", x"10", x"00", x"EE", x"0E", -- 0x17C0,
      x"4E", x"04", x"00", x"00", x"00", x"09", x"00", x"00", -- 0x17C8,
      x"00", x"00", x"00", x"00", x"00", x"00", x"EE", x"0E", -- 0x17D0,
      x"AA", x"0A", x"00", x"00", x"22", x"02", x"EE", x"0E", -- 0x17D8,
      x"EE", x"0E", x"EE", x"0E", x"EE", x"0E", x"00", x"00", -- 0x17E0,
      x"44", x"04", x"EE", x"0E", x"AA", x"0A", x"30", x"31", -- 0x17E8,
      x"32", x"33", x"34", x"35", x"36", x"37", x"38", x"39", -- 0x17F0,
      x"41", x"42", x"43", x"44", x"45", x"46", x"21", x"00", -- 0x17F8,
      x"02", x"E5", x"AF", x"F5", x"33", x"26", x"18", x"E5", -- 0x1800,
      x"CD", x"46", x"37", x"F1", x"F1", x"33", x"C9", x"21", -- 0x1808,
      x"C0", x"03", x"E5", x"3E", x"20", x"F5", x"33", x"21", -- 0x1810,
      x"00", x"00", x"E5", x"CD", x"46", x"37", x"F1", x"F1", -- 0x1818,
      x"33", x"C9", x"21", x"78", x"00", x"E5", x"3E", x"20", -- 0x1820,
      x"F5", x"33", x"21", x"48", x"03", x"E5", x"CD", x"46", -- 0x1828,
      x"37", x"F1", x"F1", x"33", x"C3", x"FE", x"17", x"FD", -- 0x1830,
      x"21", x"04", x"00", x"FD", x"39", x"FD", x"34", x"00", -- 0x1838,
      x"FD", x"4E", x"00", x"FD", x"2B", x"FD", x"2B", x"FD", -- 0x1840,
      x"5E", x"00", x"FD", x"56", x"01", x"1A", x"47", x"EE", -- 0x1848,
      x"80", x"D6", x"A0", x"38", x"12", x"0D", x"28", x"0F", -- 0x1850,
      x"78", x"D3", x"BE", x"13", x"1A", x"D6", x"2E", x"20", -- 0x1858,
      x"EC", x"3A", x"4F", x"73", x"B7", x"20", x"E6", x"79", -- 0x1860,
      x"B7", x"C8", x"0D", x"C8", x"3E", x"20", x"D3", x"BE", -- 0x1868,
      x"18", x"F8", x"CD", x"13", x"3F", x"3B", x"DD", x"36", -- 0x1870,
      x"FF", x"7E", x"DD", x"5E", x"06", x"DD", x"56", x"07", -- 0x1878,
      x"DD", x"4E", x"04", x"DD", x"46", x"05", x"1A", x"6F", -- 0x1880,
      x"B7", x"28", x"10", x"DD", x"66", x"FF", x"DD", x"35", -- 0x1888,
      x"FF", x"7C", x"B7", x"28", x"06", x"7D", x"13", x"02", -- 0x1890,
      x"03", x"18", x"EB", x"AF", x"02", x"33", x"DD", x"E1", -- 0x1898,
      x"C9", x"CD", x"B1", x"05", x"3A", x"39", x"72", x"3C", -- 0x18A0,
      x"20", x"F7", x"C9", x"CD", x"B1", x"05", x"3A", x"39", -- 0x18A8,
      x"72", x"D6", x"12", x"20", x"F6", x"C9", x"CD", x"8C", -- 0x18B0,
      x"2F", x"4D", x"21", x"02", x"00", x"39", x"7E", x"E6", -- 0x18B8,
      x"BF", x"D3", x"BF", x"3E", x"81", x"D3", x"BF", x"C5", -- 0x18C0,
      x"CD", x"B1", x"05", x"C1", x"3A", x"39", x"72", x"3C", -- 0x18C8,
      x"20", x"15", x"3A", x"3A", x"72", x"B7", x"20", x"0F", -- 0x18D0,
      x"3A", x"3B", x"72", x"B7", x"20", x"09", x"C5", x"CD", -- 0x18D8,
      x"8C", x"2F", x"7D", x"C1", x"91", x"28", x"E0", x"21", -- 0x18E0,
      x"02", x"00", x"39", x"7E", x"D3", x"BF", x"3E", x"81", -- 0x18E8,
      x"D3", x"BF", x"C9", x"CD", x"13", x"3F", x"CD", x"22", -- 0x18F0,
      x"18", x"DD", x"6E", x"04", x"DD", x"66", x"05", x"E5", -- 0x18F8,
      x"AF", x"F5", x"33", x"CD", x"38", x"08", x"33", x"21", -- 0x1900,
      x"67", x"19", x"E3", x"3E", x"01", x"F5", x"33", x"CD", -- 0x1908,
      x"38", x"08", x"F1", x"33", x"DD", x"4E", x"06", x"CB", -- 0x1910,
      x"39", x"CB", x"39", x"CB", x"39", x"CB", x"39", x"3A", -- 0x1918,
      x"4E", x"73", x"B7", x"28", x"15", x"3E", x"1E", x"D3", -- 0x1920,
      x"BF", x"AF", x"F6", x"40", x"D3", x"BF", x"79", x"D3", -- 0x1928,
      x"BE", x"DD", x"7E", x"06", x"E6", x"0F", x"D3", x"BE", -- 0x1930,
      x"18", x"1F", x"3E", x"26", x"D3", x"BF", x"AF", x"F6", -- 0x1938,
      x"40", x"D3", x"BF", x"11", x"EE", x"17", x"69", x"26", -- 0x1940,
      x"00", x"19", x"7E", x"D3", x"BE", x"DD", x"7E", x"06", -- 0x1948,
      x"E6", x"0F", x"26", x"00", x"6F", x"19", x"7E", x"D3", -- 0x1950,
      x"BE", x"CD", x"A1", x"18", x"CD", x"AB", x"18", x"CD", -- 0x1958,
      x"FE", x"17", x"DD", x"E1", x"C3", x"A1", x"18", x"50", -- 0x1960,
      x"72", x"65", x"73", x"73", x"20", x"66", x"69", x"72", -- 0x1968,
      x"65", x"2E", x"2E", x"2E", x"00", x"CD", x"13", x"3F", -- 0x1970,
      x"F5", x"DD", x"4E", x"04", x"DD", x"46", x"05", x"DD", -- 0x1978,
      x"7E", x"06", x"DD", x"77", x"FE", x"DD", x"7E", x"07", -- 0x1980,
      x"DD", x"77", x"FF", x"0A", x"5F", x"E1", x"E5", x"56", -- 0x1988,
      x"CB", x"73", x"28", x"04", x"CB", x"AB", x"18", x"07", -- 0x1990,
      x"7B", x"D6", x"5F", x"20", x"02", x"1E", x"20", x"CB", -- 0x1998,
      x"72", x"28", x"04", x"CB", x"AA", x"18", x"07", x"7A", -- 0x19A0,
      x"D6", x"5F", x"20", x"02", x"16", x"20", x"7B", x"BA", -- 0x19A8,
      x"20", x"0E", x"B7", x"28", x"0B", x"03", x"DD", x"34", -- 0x19B0,
      x"FE", x"20", x"D0", x"DD", x"34", x"FF", x"18", x"CB", -- 0x19B8,
      x"7B", x"92", x"6F", x"F1", x"DD", x"E1", x"C9", x"CD", -- 0x19C0,
      x"13", x"3F", x"F5", x"F5", x"21", x"00", x"80", x"22", -- 0x19C8,
      x"48", x"73", x"21", x"C3", x"66", x"E5", x"21", x"08", -- 0x19D0,
      x"71", x"E5", x"CD", x"9C", x"2F", x"F1", x"F1", x"7D", -- 0x19D8,
      x"B7", x"C2", x"4B", x"1B", x"21", x"C3", x"66", x"E5", -- 0x19E0,
      x"21", x"C3", x"68", x"E5", x"CD", x"72", x"18", x"F1", -- 0x19E8,
      x"21", x"C3", x"68", x"E3", x"3E", x"01", x"F5", x"33", -- 0x19F0,
      x"CD", x"38", x"08", x"F1", x"33", x"3A", x"C4", x"66", -- 0x19F8,
      x"B7", x"28", x"33", x"2A", x"48", x"73", x"DD", x"75", -- 0x1A00,
      x"FE", x"DD", x"74", x"FF", x"21", x"80", x"00", x"E5", -- 0x1A08,
      x"2E", x"00", x"E5", x"DD", x"6E", x"FE", x"DD", x"66", -- 0x1A10,
      x"FF", x"E5", x"CD", x"D1", x"00", x"F1", x"F1", x"F1", -- 0x1A18,
      x"2A", x"48", x"73", x"36", x"2E", x"2A", x"48", x"73", -- 0x1A20,
      x"23", x"36", x"2E", x"21", x"48", x"73", x"7E", x"C6", -- 0x1A28,
      x"80", x"77", x"30", x"02", x"23", x"34", x"11", x"34", -- 0x1A30,
      x"71", x"01", x"08", x"71", x"D5", x"C5", x"CD", x"F4", -- 0x1A38,
      x"4A", x"F1", x"F1", x"7D", x"B7", x"C2", x"3E", x"1B", -- 0x1A40,
      x"CD", x"8C", x"2F", x"7D", x"D6", x"02", x"20", x"0B", -- 0x1A48,
      x"01", x"08", x"71", x"C5", x"CD", x"55", x"46", x"F1", -- 0x1A50,
      x"C3", x"4B", x"1B", x"3A", x"39", x"71", x"FE", x"2E", -- 0x1A58,
      x"28", x"D4", x"B7", x"CA", x"3E", x"1B", x"3A", x"4D", -- 0x1A60,
      x"73", x"B7", x"28", x"3D", x"3A", x"38", x"71", x"CB", -- 0x1A68,
      x"67", x"28", x"36", x"21", x"B6", x"17", x"E5", x"21", -- 0x1A70,
      x"39", x"71", x"E5", x"CD", x"75", x"19", x"F1", x"F1", -- 0x1A78,
      x"7D", x"B7", x"20", x"25", x"21", x"08", x"71", x"E5", -- 0x1A80,
      x"CD", x"55", x"46", x"F1", x"21", x"BD", x"17", x"4E", -- 0x1A88,
      x"06", x"00", x"C5", x"21", x"B6", x"17", x"E5", x"21", -- 0x1A90,
      x"C4", x"66", x"E5", x"CD", x"AE", x"00", x"F1", x"F1", -- 0x1A98,
      x"F1", x"21", x"4D", x"73", x"36", x"00", x"C3", x"CC", -- 0x1AA0,
      x"19", x"21", x"39", x"71", x"E5", x"2A", x"48", x"73", -- 0x1AA8,
      x"E5", x"CD", x"72", x"18", x"F1", x"F1", x"21", x"38", -- 0x1AB0,
      x"71", x"5E", x"FD", x"21", x"48", x"73", x"FD", x"7E", -- 0x1AB8,
      x"00", x"C6", x"7F", x"4F", x"FD", x"7E", x"01", x"CE", -- 0x1AC0,
      x"00", x"47", x"CB", x"63", x"28", x"04", x"AF", x"02", -- 0x1AC8,
      x"18", x"33", x"C5", x"11", x"34", x"71", x"21", x"02", -- 0x1AD0,
      x"00", x"39", x"EB", x"01", x"04", x"00", x"ED", x"B0", -- 0x1AD8,
      x"C1", x"DD", x"5E", x"FD", x"DD", x"56", x"FE", x"DD", -- 0x1AE0,
      x"6E", x"FF", x"3E", x"06", x"CB", x"3D", x"CB", x"1A", -- 0x1AE8,
      x"CB", x"1B", x"3D", x"20", x"F7", x"DD", x"7E", x"FC", -- 0x1AF0,
      x"B7", x"20", x"07", x"DD", x"7E", x"FD", x"E6", x"3F", -- 0x1AF8,
      x"28", x"01", x"1C", x"7B", x"02", x"21", x"48", x"73", -- 0x1B00,
      x"7E", x"C6", x"80", x"77", x"30", x"02", x"23", x"34", -- 0x1B08,
      x"FD", x"21", x"48", x"73", x"FD", x"7E", x"00", x"D6", -- 0x1B10,
      x"80", x"FD", x"7E", x"01", x"DE", x"FF", x"DA", x"36", -- 0x1B18,
      x"1A", x"ED", x"4B", x"48", x"73", x"59", x"78", x"C6", -- 0x1B20,
      x"80", x"57", x"06", x"07", x"CB", x"3A", x"CB", x"1B", -- 0x1B28,
      x"10", x"FA", x"7B", x"F5", x"33", x"21", x"50", x"1B", -- 0x1B30,
      x"E5", x"CD", x"F3", x"18", x"F1", x"33", x"21", x"08", -- 0x1B38,
      x"71", x"E5", x"CD", x"55", x"46", x"F1", x"21", x"4D", -- 0x1B40,
      x"73", x"36", x"00", x"DD", x"F9", x"DD", x"E1", x"C9", -- 0x1B48,
      x"4D", x"61", x"78", x"20", x"64", x"69", x"72", x"65", -- 0x1B50,
      x"63", x"74", x"6F", x"72", x"79", x"20", x"63", x"6F", -- 0x1B58,
      x"75", x"6E", x"74", x"20", x"72", x"65", x"61", x"63", -- 0x1B60,
      x"68", x"65", x"64", x"00", x"CD", x"B1", x"05", x"3A", -- 0x1B68,
      x"3A", x"72", x"B7", x"20", x"0C", x"3A", x"3B", x"72", -- 0x1B70,
      x"B7", x"20", x"06", x"21", x"C3", x"6C", x"36", x"2D", -- 0x1B78,
      x"C9", x"FD", x"21", x"C3", x"6C", x"FD", x"35", x"00", -- 0x1B80,
      x"FD", x"7E", x"00", x"B7", x"20", x"05", x"FD", x"36", -- 0x1B88,
      x"00", x"05", x"C9", x"3E", x"01", x"F5", x"33", x"CD", -- 0x1B90,
      x"7A", x"02", x"33", x"18", x"CF", x"CD", x"13", x"3F", -- 0x1B98,
      x"21", x"F7", x"FF", x"39", x"F9", x"3A", x"4B", x"73", -- 0x1BA0,
      x"DD", x"77", x"FB", x"DD", x"36", x"FC", x"00", x"DD", -- 0x1BA8,
      x"36", x"FD", x"10", x"AF", x"DD", x"77", x"FE", x"DD", -- 0x1BB0,
      x"77", x"FF", x"21", x"4B", x"73", x"4E", x"06", x"00", -- 0x1BB8,
      x"21", x"18", x"00", x"09", x"DD", x"7E", x"FB", x"DD", -- 0x1BC0,
      x"77", x"F7", x"AF", x"DD", x"77", x"F8", x"DD", x"7E", -- 0x1BC8,
      x"F7", x"95", x"DD", x"7E", x"F8", x"9C", x"E2", x"DB", -- 0x1BD0,
      x"1B", x"EE", x"80", x"F2", x"DD", x"1C", x"DD", x"7E", -- 0x1BD8,
      x"FB", x"E6", x"01", x"DD", x"77", x"F9", x"DD", x"36", -- 0x1BE0,
      x"FA", x"00", x"3E", x"00", x"DD", x"B6", x"F9", x"28", -- 0x1BE8,
      x"17", x"21", x"28", x"00", x"E5", x"3E", x"43", x"F5", -- 0x1BF0,
      x"33", x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"E5", -- 0x1BF8,
      x"CD", x"46", x"37", x"F1", x"F1", x"33", x"18", x"15", -- 0x1C00,
      x"21", x"28", x"00", x"E5", x"3E", x"42", x"F5", x"33", -- 0x1C08,
      x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"E5", x"CD", -- 0x1C10,
      x"46", x"37", x"F1", x"F1", x"33", x"DD", x"46", x"FF", -- 0x1C18,
      x"DD", x"4E", x"FE", x"CB", x"F0", x"21", x"4A", x"73", -- 0x1C20,
      x"DD", x"7E", x"FB", x"96", x"38", x"2D", x"79", x"D3", -- 0x1C28,
      x"BF", x"78", x"D3", x"BF", x"3E", x"28", x"F5", x"33", -- 0x1C30,
      x"21", x"E2", x"1C", x"E5", x"CD", x"37", x"18", x"F1", -- 0x1C38,
      x"33", x"DD", x"7E", x"FB", x"3C", x"20", x"76", x"DD", -- 0x1C40,
      x"35", x"FB", x"DD", x"7E", x"FE", x"D6", x"98", x"20", -- 0x1C48,
      x"6C", x"DD", x"7E", x"FF", x"D6", x"03", x"CA", x"DD", -- 0x1C50,
      x"1C", x"18", x"62", x"E1", x"E5", x"29", x"11", x"C3", -- 0x1C58,
      x"6A", x"19", x"5E", x"23", x"56", x"6B", x"62", x"C5", -- 0x1C60,
      x"01", x"7F", x"00", x"09", x"C1", x"7E", x"B7", x"20", -- 0x1C68,
      x"3C", x"DD", x"7E", x"FA", x"DD", x"B6", x"F9", x"28", -- 0x1C70,
      x"1B", x"C5", x"D5", x"21", x"28", x"00", x"E5", x"3E", -- 0x1C78,
      x"53", x"F5", x"33", x"DD", x"6E", x"FC", x"DD", x"66", -- 0x1C80,
      x"FD", x"E5", x"CD", x"46", x"37", x"F1", x"F1", x"33", -- 0x1C88,
      x"D1", x"C1", x"18", x"19", x"C5", x"D5", x"21", x"28", -- 0x1C90,
      x"00", x"E5", x"3E", x"52", x"F5", x"33", x"DD", x"6E", -- 0x1C98,
      x"FC", x"DD", x"66", x"FD", x"E5", x"CD", x"46", x"37", -- 0x1CA0,
      x"F1", x"F1", x"33", x"D1", x"C1", x"79", x"D3", x"BF", -- 0x1CA8,
      x"78", x"D3", x"BF", x"3E", x"28", x"F5", x"33", x"D5", -- 0x1CB0,
      x"CD", x"37", x"18", x"F1", x"33", x"DD", x"7E", x"FC", -- 0x1CB8,
      x"C6", x"28", x"DD", x"77", x"FC", x"30", x"03", x"DD", -- 0x1CC0,
      x"34", x"FD", x"DD", x"7E", x"FE", x"C6", x"28", x"DD", -- 0x1CC8,
      x"77", x"FE", x"30", x"03", x"DD", x"34", x"FF", x"DD", -- 0x1CD0,
      x"34", x"FB", x"C3", x"BA", x"1B", x"DD", x"F9", x"DD", -- 0x1CD8,
      x"E1", x"C9", x"00", x"CD", x"13", x"3F", x"F5", x"F5", -- 0x1CE0,
      x"21", x"4A", x"73", x"36", x"00", x"DD", x"36", x"FE", -- 0x1CE8,
      x"00", x"DD", x"36", x"FF", x"80", x"21", x"48", x"73", -- 0x1CF0,
      x"DD", x"7E", x"FE", x"96", x"DD", x"7E", x"FF", x"23", -- 0x1CF8,
      x"9E", x"D2", x"EF", x"1D", x"C1", x"E1", x"E5", x"C5", -- 0x1D00,
      x"11", x"7F", x"00", x"19", x"7E", x"B7", x"20", x"35", -- 0x1D08,
      x"4F", x"21", x"4A", x"73", x"79", x"96", x"30", x"66", -- 0x1D10,
      x"69", x"26", x"00", x"29", x"11", x"C3", x"6A", x"19", -- 0x1D18,
      x"5E", x"23", x"56", x"6B", x"62", x"C5", x"01", x"7F", -- 0x1D20,
      x"00", x"09", x"C1", x"7E", x"B7", x"20", x"4F", x"C5", -- 0x1D28,
      x"D5", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"E5", -- 0x1D30,
      x"CD", x"75", x"19", x"F1", x"F1", x"C1", x"CB", x"7D", -- 0x1D38,
      x"20", x"3C", x"0C", x"18", x"CC", x"21", x"4A", x"73", -- 0x1D40,
      x"4E", x"0D", x"41", x"78", x"3C", x"28", x"2F", x"68", -- 0x1D48,
      x"26", x"00", x"29", x"11", x"C3", x"6A", x"19", x"5E", -- 0x1D50,
      x"23", x"56", x"6B", x"62", x"C5", x"01", x"7F", x"00", -- 0x1D58,
      x"09", x"C1", x"7E", x"0C", x"B7", x"28", x"17", x"C5", -- 0x1D60,
      x"D5", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"E5", -- 0x1D68,
      x"CD", x"75", x"19", x"F1", x"F1", x"C1", x"CB", x"7D", -- 0x1D70,
      x"28", x"04", x"05", x"48", x"18", x"CD", x"59", x"16", -- 0x1D78,
      x"00", x"DD", x"73", x"FC", x"DD", x"72", x"FD", x"DD", -- 0x1D80,
      x"CB", x"FC", x"26", x"DD", x"CB", x"FD", x"16", x"21", -- 0x1D88,
      x"4A", x"73", x"79", x"96", x"30", x"2F", x"FD", x"21", -- 0x1D90,
      x"4A", x"73", x"FD", x"6E", x"00", x"26", x"00", x"BF", -- 0x1D98,
      x"ED", x"52", x"29", x"3E", x"C3", x"DD", x"86", x"FC", -- 0x1DA0,
      x"4F", x"3E", x"6A", x"DD", x"8E", x"FD", x"47", x"13", -- 0x1DA8,
      x"CB", x"23", x"CB", x"12", x"7B", x"C6", x"C3", x"5F", -- 0x1DB0,
      x"7A", x"CE", x"6A", x"57", x"E5", x"C5", x"D5", x"CD", -- 0x1DB8,
      x"0B", x"01", x"F1", x"F1", x"F1", x"DD", x"7E", x"FC", -- 0x1DC0,
      x"C6", x"C3", x"4F", x"DD", x"7E", x"FD", x"CE", x"6A", -- 0x1DC8,
      x"47", x"DD", x"7E", x"FE", x"02", x"03", x"DD", x"7E", -- 0x1DD0,
      x"FF", x"02", x"21", x"4A", x"73", x"34", x"DD", x"7E", -- 0x1DD8,
      x"FE", x"C6", x"80", x"DD", x"77", x"FE", x"D2", x"F5", -- 0x1DE0,
      x"1C", x"DD", x"34", x"FF", x"C3", x"F5", x"1C", x"DD", -- 0x1DE8,
      x"F9", x"DD", x"E1", x"C9", x"3B", x"CD", x"FE", x"17", -- 0x1DF0,
      x"21", x"77", x"1E", x"E5", x"21", x"40", x"18", x"E5", -- 0x1DF8,
      x"CD", x"35", x"06", x"F1", x"21", x"90", x"1E", x"E3", -- 0x1E00,
      x"21", x"18", x"18", x"E5", x"CD", x"35", x"06", x"F1", -- 0x1E08,
      x"F1", x"01", x"18", x"15", x"AF", x"FD", x"21", x"00", -- 0x1E10,
      x"00", x"FD", x"39", x"FD", x"77", x"00", x"21", x"00", -- 0x1E18,
      x"00", x"39", x"7E", x"D6", x"02", x"30", x"4E", x"C5", -- 0x1E20,
      x"3E", x"02", x"F5", x"33", x"CD", x"7A", x"02", x"33", -- 0x1E28,
      x"C1", x"59", x"50", x"1B", x"4B", x"7A", x"47", x"B3", -- 0x1E30,
      x"20", x"15", x"3E", x"E2", x"F5", x"33", x"CD", x"B6", -- 0x1E38,
      x"18", x"33", x"01", x"18", x"15", x"AF", x"FD", x"21", -- 0x1E40,
      x"00", x"00", x"FD", x"39", x"FD", x"77", x"00", x"C5", -- 0x1E48,
      x"CD", x"8C", x"2F", x"7D", x"C1", x"D6", x"02", x"20", -- 0x1E50,
      x"0C", x"AF", x"FD", x"21", x"00", x"00", x"FD", x"39", -- 0x1E58,
      x"FD", x"77", x"00", x"18", x"09", x"FD", x"21", x"00", -- 0x1E60,
      x"00", x"FD", x"39", x"FD", x"34", x"00", x"C5", x"CD", -- 0x1E68,
      x"B1", x"05", x"C1", x"18", x"A9", x"33", x"C9", x"49", -- 0x1E70,
      x"6E", x"73", x"65", x"72", x"74", x"20", x"53", x"44", -- 0x1E78,
      x"20", x"6F", x"72", x"20", x"74", x"75", x"72", x"6E", -- 0x1E80,
      x"20", x"73", x"79", x"73", x"74", x"65", x"6D", x"00", -- 0x1E88,
      x"6F", x"66", x"66", x"20", x"62", x"65", x"66", x"6F", -- 0x1E90,
      x"72", x"65", x"20", x"69", x"6E", x"73", x"65", x"72", -- 0x1E98,
      x"74", x"69", x"6E", x"67", x"20", x"63", x"61", x"72", -- 0x1EA0,
      x"74", x"72", x"69", x"64", x"67", x"65", x"00", x"CD", -- 0x1EA8,
      x"13", x"3F", x"F5", x"F5", x"F5", x"CD", x"22", x"18", -- 0x1EB0,
      x"21", x"60", x"1F", x"E5", x"AF", x"F5", x"33", x"CD", -- 0x1EB8,
      x"38", x"08", x"F1", x"33", x"11", x"00", x"82", x"21", -- 0x1EC0,
      x"00", x"00", x"39", x"4B", x"42", x"D5", x"E5", x"21", -- 0x1EC8,
      x"00", x"02", x"E5", x"C5", x"21", x"EC", x"6E", x"E5", -- 0x1ED0,
      x"CD", x"DC", x"29", x"F1", x"F1", x"F1", x"F1", x"7D", -- 0x1ED8,
      x"D1", x"47", x"B7", x"28", x"14", x"C5", x"21", x"EC", -- 0x1EE0,
      x"6E", x"E5", x"CD", x"7B", x"46", x"33", x"21", x"70", -- 0x1EE8,
      x"1F", x"E3", x"CD", x"F3", x"18", x"F1", x"33", x"18", -- 0x1EF0,
      x"62", x"DD", x"7E", x"FB", x"D6", x"02", x"38", x"4C", -- 0x1EF8,
      x"21", x"00", x"02", x"19", x"EB", x"7A", x"D6", x"80", -- 0x1F00,
      x"30", x"BD", x"11", x"FC", x"6E", x"21", x"02", x"00", -- 0x1F08,
      x"39", x"EB", x"01", x"04", x"00", x"ED", x"B0", x"ED", -- 0x1F10,
      x"4B", x"F6", x"6E", x"ED", x"5B", x"F8", x"6E", x"DD", -- 0x1F18,
      x"7E", x"FC", x"91", x"20", x"11", x"DD", x"7E", x"FD", -- 0x1F20,
      x"90", x"20", x"0B", x"DD", x"6E", x"FE", x"DD", x"66", -- 0x1F28,
      x"FF", x"BF", x"ED", x"52", x"28", x"16", x"21", x"EC", -- 0x1F30,
      x"6E", x"E5", x"CD", x"7B", x"46", x"26", x"01", x"E3", -- 0x1F38,
      x"33", x"21", x"87", x"1F", x"E5", x"CD", x"F3", x"18", -- 0x1F40,
      x"F1", x"33", x"18", x"0F", x"21", x"EC", x"6E", x"E5", -- 0x1F48,
      x"CD", x"7B", x"46", x"F1", x"3E", x"31", x"D3", x"55", -- 0x1F50,
      x"CD", x"C2", x"08", x"DD", x"F9", x"DD", x"E1", x"C9", -- 0x1F58,
      x"72", x"65", x"61", x"64", x"69", x"6E", x"67", x"20", -- 0x1F60,
      x"63", x"61", x"72", x"74", x"2E", x"2E", x"2E", x"00", -- 0x1F68,
      x"43", x"61", x"72", x"74", x"72", x"69", x"64", x"67", -- 0x1F70,
      x"65", x"20", x"6C", x"6F", x"61", x"64", x"20", x"66", -- 0x1F78,
      x"61", x"69", x"6C", x"65", x"64", x"2E", x"00", x"55", -- 0x1F80,
      x"6E", x"72", x"65", x"63", x"6F", x"67", x"6E", x"69", -- 0x1F88,
      x"7A", x"65", x"64", x"20", x"3E", x"33", x"32", x"6B", -- 0x1F90,
      x"20", x"43", x"61", x"72", x"74", x"00", x"CD", x"13", -- 0x1F98,
      x"3F", x"01", x"80", x"00", x"79", x"B0", x"28", x"36", -- 0x1FA0,
      x"DD", x"7E", x"04", x"D3", x"54", x"58", x"51", x"C5", -- 0x1FA8,
      x"D5", x"21", x"00", x"02", x"E5", x"D5", x"21", x"C3", -- 0x1FB0,
      x"68", x"E5", x"CD", x"AE", x"00", x"F1", x"F1", x"F1", -- 0x1FB8,
      x"D1", x"C1", x"DD", x"7E", x"05", x"D3", x"54", x"C5", -- 0x1FC0,
      x"21", x"00", x"02", x"E5", x"21", x"C3", x"68", x"E5", -- 0x1FC8,
      x"D5", x"CD", x"AE", x"00", x"F1", x"F1", x"F1", x"C1", -- 0x1FD0,
      x"79", x"C6", x"02", x"4F", x"18", x"C6", x"DD", x"E1", -- 0x1FD8,
      x"C9", x"CD", x"13", x"3F", x"21", x"F6", x"FF", x"39", -- 0x1FE0,
      x"F9", x"CD", x"22", x"18", x"21", x"9B", x"21", x"E5", -- 0x1FE8,
      x"AF", x"F5", x"33", x"CD", x"38", x"08", x"F1", x"33", -- 0x1FF0,
      x"11", x"00", x"00", x"01", x"00", x"00", x"DD", x"7E", -- 0x1FF8,
      x"04", x"D6", x"20", x"20", x"0E", x"11", x"00", x"80", -- 0x2000,
      x"01", x"00", x"00", x"DD", x"7E", x"04", x"C6", x"FE", -- 0x2008,
      x"DD", x"77", x"04", x"DD", x"6E", x"04", x"26", x"00", -- 0x2010,
      x"2B", x"CB", x"2C", x"CB", x"1D", x"3E", x"0F", x"95", -- 0x2018,
      x"DD", x"77", x"FC", x"D3", x"54", x"DD", x"7E", x"04", -- 0x2020,
      x"0F", x"30", x"05", x"21", x"00", x"40", x"18", x"03", -- 0x2028,
      x"21", x"00", x"00", x"DD", x"75", x"FD", x"7C", x"C6", -- 0x2030,
      x"80", x"DD", x"77", x"FE", x"C5", x"D5", x"21", x"EC", -- 0x2038,
      x"6E", x"E5", x"CD", x"46", x"3F", x"F1", x"F1", x"F1", -- 0x2040,
      x"7D", x"B7", x"28", x"1A", x"21", x"EC", x"6E", x"E5", -- 0x2048,
      x"CD", x"7B", x"46", x"26", x"02", x"E3", x"33", x"21", -- 0x2050,
      x"AF", x"21", x"E5", x"CD", x"F3", x"18", x"F1", x"33", -- 0x2058,
      x"DD", x"6E", x"FC", x"C3", x"96", x"21", x"DD", x"7E", -- 0x2060,
      x"FC", x"DD", x"77", x"FF", x"21", x"04", x"00", x"39", -- 0x2068,
      x"DD", x"4E", x"FD", x"DD", x"46", x"FE", x"E5", x"21", -- 0x2070,
      x"00", x"02", x"E5", x"C5", x"21", x"EC", x"6E", x"E5", -- 0x2078,
      x"CD", x"DC", x"29", x"F1", x"F1", x"F1", x"F1", x"7D", -- 0x2080,
      x"47", x"B7", x"28", x"18", x"C5", x"21", x"EC", x"6E", -- 0x2088,
      x"E5", x"CD", x"7B", x"46", x"33", x"21", x"C4", x"21", -- 0x2090,
      x"E3", x"CD", x"F3", x"18", x"F1", x"33", x"DD", x"6E", -- 0x2098,
      x"FC", x"C3", x"96", x"21", x"DD", x"7E", x"FB", x"D6", -- 0x20A0,
      x"02", x"38", x"78", x"DD", x"7E", x"FD", x"DD", x"77", -- 0x20A8,
      x"FD", x"DD", x"7E", x"FE", x"C6", x"02", x"DD", x"77", -- 0x20B0,
      x"FE", x"D6", x"80", x"30", x"AF", x"DD", x"34", x"FF", -- 0x20B8,
      x"DD", x"7E", x"FF", x"DD", x"77", x"FC", x"3E", x"0F", -- 0x20C0,
      x"DD", x"96", x"FF", x"30", x"46", x"11", x"FC", x"6E", -- 0x20C8,
      x"21", x"00", x"00", x"39", x"EB", x"01", x"04", x"00", -- 0x20D0,
      x"ED", x"B0", x"ED", x"4B", x"F6", x"6E", x"ED", x"5B", -- 0x20D8,
      x"F8", x"6E", x"DD", x"7E", x"F6", x"91", x"20", x"11", -- 0x20E0,
      x"DD", x"7E", x"F7", x"90", x"20", x"0B", x"DD", x"6E", -- 0x20E8,
      x"F8", x"DD", x"66", x"F9", x"BF", x"ED", x"52", x"28", -- 0x20F0,
      x"2A", x"21", x"EC", x"6E", x"E5", x"CD", x"7B", x"46", -- 0x20F8,
      x"F1", x"AF", x"F5", x"33", x"21", x"DB", x"21", x"E5", -- 0x2100,
      x"CD", x"F3", x"18", x"F1", x"33", x"DD", x"6E", x"FF", -- 0x2108,
      x"C3", x"96", x"21", x"DD", x"36", x"FD", x"00", x"DD", -- 0x2110,
      x"36", x"FE", x"80", x"DD", x"7E", x"FF", x"D3", x"54", -- 0x2118,
      x"C3", x"6C", x"20", x"21", x"EC", x"6E", x"E5", x"CD", -- 0x2120,
      x"7B", x"46", x"F1", x"DD", x"7E", x"04", x"D6", x"02", -- 0x2128,
      x"28", x"1E", x"DD", x"7E", x"04", x"D6", x"04", x"28", -- 0x2130,
      x"1D", x"DD", x"7E", x"04", x"D6", x"08", x"28", x"1C", -- 0x2138,
      x"DD", x"7E", x"04", x"D6", x"10", x"28", x"1B", x"DD", -- 0x2140,
      x"7E", x"04", x"D6", x"1E", x"28", x"1A", x"18", x"1E", -- 0x2148,
      x"3E", x"01", x"D3", x"59", x"18", x"33", x"3E", x"03", -- 0x2150,
      x"D3", x"59", x"18", x"2D", x"3E", x"07", x"D3", x"59", -- 0x2158,
      x"18", x"27", x"3E", x"0F", x"D3", x"59", x"18", x"21", -- 0x2160,
      x"3E", x"1F", x"D3", x"59", x"18", x"1B", x"21", x"EC", -- 0x2168,
      x"6E", x"E5", x"CD", x"7B", x"46", x"F1", x"DD", x"7E", -- 0x2170,
      x"04", x"F5", x"33", x"21", x"F2", x"21", x"E5", x"CD", -- 0x2178,
      x"F3", x"18", x"F1", x"33", x"DD", x"6E", x"FC", x"18", -- 0x2180,
      x"0D", x"3E", x"11", x"D3", x"55", x"3E", x"01", x"D3", -- 0x2188,
      x"54", x"CD", x"C2", x"08", x"2E", x"00", x"DD", x"F9", -- 0x2190,
      x"DD", x"E1", x"C9", x"72", x"65", x"61", x"64", x"69", -- 0x2198,
      x"6E", x"67", x"20", x"6D", x"65", x"67", x"61", x"63", -- 0x21A0,
      x"61", x"72", x"74", x"2E", x"2E", x"2E", x"00", x"46", -- 0x21A8,
      x"61", x"69", x"6C", x"65", x"64", x"20", x"74", x"6F", -- 0x21B0,
      x"20", x"73", x"65", x"65", x"6B", x"20", x"66", x"69", -- 0x21B8,
      x"6C", x"65", x"2E", x"00", x"43", x"61", x"72", x"74", -- 0x21C0,
      x"72", x"69", x"64", x"67", x"65", x"20", x"6C", x"6F", -- 0x21C8,
      x"61", x"64", x"20", x"66", x"61", x"69", x"6C", x"65", -- 0x21D0,
      x"64", x"2E", x"00", x"4D", x"65", x"67", x"61", x"63", -- 0x21D8,
      x"61", x"72", x"74", x"20", x"52", x"4F", x"4D", x"20", -- 0x21E0,
      x"74", x"6F", x"6F", x"20", x"6C", x"61", x"72", x"67", -- 0x21E8,
      x"65", x"00", x"4D", x"65", x"67", x"61", x"63", x"61", -- 0x21F0,
      x"72", x"74", x"20", x"69", x"6D", x"61", x"67", x"65", -- 0x21F8,
      x"73", x"20", x"6D", x"75", x"73", x"74", x"20", x"62", -- 0x2200,
      x"65", x"20", x"70", x"61", x"64", x"64", x"65", x"64", -- 0x2208,
      x"00", x"21", x"4A", x"73", x"4E", x"06", x"00", x"0B", -- 0x2210,
      x"21", x"4C", x"73", x"5E", x"16", x"00", x"79", x"93", -- 0x2218,
      x"78", x"9A", x"E2", x"27", x"22", x"EE", x"80", x"F2", -- 0x2220,
      x"33", x"22", x"3A", x"4A", x"73", x"21", x"4C", x"73", -- 0x2228,
      x"C6", x"FF", x"77", x"21", x"4C", x"73", x"4E", x"06", -- 0x2230,
      x"00", x"21", x"4B", x"73", x"5E", x"16", x"00", x"79", -- 0x2238,
      x"93", x"4F", x"78", x"9A", x"47", x"69", x"60", x"29", -- 0x2240,
      x"29", x"09", x"29", x"29", x"29", x"4D", x"7C", x"C6", -- 0x2248,
      x"10", x"47", x"C5", x"C5", x"CD", x"DC", x"33", x"F1", -- 0x2250,
      x"7D", x"C1", x"E6", x"F0", x"F6", x"07", x"57", x"21", -- 0x2258,
      x"28", x"00", x"E5", x"D5", x"33", x"C5", x"CD", x"46", -- 0x2260,
      x"37", x"F1", x"F1", x"33", x"C9", x"21", x"4C", x"73", -- 0x2268,
      x"4E", x"06", x"00", x"21", x"4B", x"73", x"5E", x"16", -- 0x2270,
      x"00", x"79", x"93", x"4F", x"78", x"9A", x"47", x"CB", -- 0x2278,
      x"41", x"1E", x"03", x"20", x"02", x"1E", x"02", x"69", -- 0x2280,
      x"60", x"29", x"29", x"09", x"29", x"29", x"29", x"4D", -- 0x2288,
      x"7C", x"C6", x"10", x"47", x"C5", x"D5", x"C5", x"CD", -- 0x2290,
      x"DC", x"33", x"F1", x"7D", x"D1", x"C1", x"E6", x"F0", -- 0x2298,
      x"B3", x"57", x"21", x"28", x"00", x"E5", x"D5", x"33", -- 0x22A0,
      x"C5", x"CD", x"46", x"37", x"F1", x"F1", x"33", x"C9", -- 0x22A8,
      x"CD", x"13", x"3F", x"F5", x"21", x"18", x"15", x"E3", -- 0x22B0,
      x"CD", x"11", x"22", x"CD", x"8C", x"2F", x"7D", x"D6", -- 0x22B8,
      x"02", x"20", x"04", x"6F", x"C3", x"27", x"24", x"3E", -- 0x22C0,
      x"01", x"F5", x"33", x"CD", x"7A", x"02", x"33", x"CD", -- 0x22C8,
      x"B1", x"05", x"3A", x"3B", x"72", x"21", x"3A", x"72", -- 0x22D0,
      x"B6", x"B7", x"CA", x"FD", x"23", x"CD", x"6D", x"22", -- 0x22D8,
      x"3A", x"3B", x"72", x"D6", x"80", x"20", x"05", x"2E", -- 0x22E0,
      x"FF", x"C3", x"27", x"24", x"3A", x"3A", x"72", x"D6", -- 0x22E8,
      x"04", x"20", x"21", x"FD", x"21", x"4C", x"73", x"FD", -- 0x22F0,
      x"7E", x"00", x"B7", x"CA", x"F0", x"23", x"FD", x"35", -- 0x22F8,
      x"00", x"21", x"4B", x"73", x"FD", x"7E", x"00", x"96", -- 0x2300,
      x"D2", x"F0", x"23", x"21", x"4B", x"73", x"35", x"2E", -- 0x2308,
      x"FF", x"C3", x"27", x"24", x"21", x"4A", x"73", x"5E", -- 0x2310,
      x"16", x"00", x"21", x"4B", x"73", x"4E", x"06", x"00", -- 0x2318,
      x"1B", x"21", x"17", x"00", x"09", x"E3", x"3A", x"3A", -- 0x2320,
      x"72", x"D6", x"FC", x"20", x"35", x"3A", x"4C", x"73", -- 0x2328,
      x"06", x"00", x"93", x"78", x"9A", x"E2", x"3A", x"23", -- 0x2330,
      x"EE", x"80", x"F2", x"F0", x"23", x"FD", x"21", x"4C", -- 0x2338,
      x"73", x"FD", x"34", x"00", x"FD", x"4E", x"00", x"06", -- 0x2340,
      x"00", x"DD", x"7E", x"FE", x"91", x"DD", x"7E", x"FF", -- 0x2348,
      x"98", x"E2", x"56", x"23", x"EE", x"80", x"F2", x"F0", -- 0x2350,
      x"23", x"21", x"4B", x"73", x"34", x"2E", x"FF", x"C3", -- 0x2358,
      x"27", x"24", x"21", x"4B", x"73", x"4E", x"21", x"4C", -- 0x2360,
      x"73", x"46", x"3A", x"3B", x"72", x"D6", x"04", x"20", -- 0x2368,
      x"45", x"FD", x"21", x"4A", x"73", x"FD", x"6E", x"00", -- 0x2370,
      x"2D", x"DD", x"7E", x"FE", x"93", x"DD", x"7E", x"FF", -- 0x2378,
      x"9A", x"E2", x"86", x"23", x"EE", x"80", x"F2", x"AD", -- 0x2380,
      x"23", x"7D", x"91", x"FE", x"18", x"30", x"0D", x"21", -- 0x2388,
      x"4B", x"73", x"86", x"77", x"3A", x"4B", x"73", x"32", -- 0x2390,
      x"4C", x"73", x"18", x"0C", x"79", x"C6", x"18", x"32", -- 0x2398,
      x"4B", x"73", x"78", x"C6", x"18", x"32", x"4C", x"73", -- 0x23A0,
      x"2E", x"FF", x"C3", x"27", x"24", x"FD", x"21", x"4C", -- 0x23A8,
      x"73", x"FD", x"75", x"00", x"18", x"3A", x"3A", x"3B", -- 0x23B0,
      x"72", x"D6", x"FC", x"20", x"33", x"FD", x"21", x"4B", -- 0x23B8,
      x"73", x"FD", x"7E", x"00", x"B7", x"28", x"24", x"FD", -- 0x23C0,
      x"7E", x"00", x"D6", x"18", x"30", x"0B", x"FD", x"36", -- 0x23C8,
      x"00", x"00", x"21", x"4C", x"73", x"36", x"00", x"18", -- 0x23D0,
      x"0E", x"21", x"4B", x"73", x"79", x"C6", x"E8", x"77", -- 0x23D8,
      x"21", x"4C", x"73", x"78", x"C6", x"E8", x"77", x"2E", -- 0x23E0,
      x"FF", x"18", x"3C", x"21", x"4C", x"73", x"36", x"00", -- 0x23E8,
      x"CD", x"11", x"22", x"CD", x"6C", x"1B", x"21", x"18", -- 0x23F0,
      x"15", x"E3", x"C3", x"BB", x"22", x"21", x"C3", x"6C", -- 0x23F8,
      x"36", x"2D", x"3A", x"39", x"72", x"D6", x"12", x"20", -- 0x2400,
      x"04", x"2E", x"01", x"18", x"1A", x"C1", x"C5", x"0B", -- 0x2408,
      x"33", x"33", x"C5", x"78", x"B1", x"C2", x"BB", x"22", -- 0x2410,
      x"3E", x"F2", x"F5", x"33", x"CD", x"B6", x"18", x"33", -- 0x2418,
      x"21", x"18", x"15", x"E3", x"C3", x"BB", x"22", x"F1", -- 0x2420,
      x"DD", x"E1", x"C9", x"01", x"50", x"73", x"FD", x"21", -- 0x2428,
      x"38", x"72", x"FD", x"6E", x"00", x"26", x"00", x"29", -- 0x2430,
      x"09", x"4E", x"23", x"46", x"3E", x"08", x"F5", x"33", -- 0x2438,
      x"C5", x"CD", x"7D", x"14", x"F1", x"33", x"C9", x"FD", -- 0x2440,
      x"21", x"38", x"72", x"FD", x"34", x"00", x"FD", x"7E", -- 0x2448,
      x"00", x"D6", x"03", x"DA", x"2B", x"24", x"FD", x"36", -- 0x2450,
      x"00", x"00", x"C3", x"2B", x"24", x"CD", x"13", x"3F", -- 0x2458,
      x"F5", x"F5", x"F5", x"CD", x"FE", x"17", x"CD", x"8C", -- 0x2460,
      x"2F", x"7D", x"D6", x"02", x"20", x"03", x"CD", x"F4", -- 0x2468,
      x"1D", x"21", x"C3", x"66", x"36", x"2F", x"21", x"C4", -- 0x2470,
      x"66", x"36", x"00", x"3E", x"01", x"F5", x"33", x"21", -- 0x2478,
      x"4D", x"28", x"E5", x"21", x"C4", x"6C", x"E5", x"CD", -- 0x2480,
      x"F2", x"31", x"F1", x"F1", x"33", x"7D", x"B7", x"28", -- 0x2488,
      x"0E", x"AF", x"F5", x"33", x"21", x"4E", x"28", x"E5", -- 0x2490,
      x"CD", x"F3", x"18", x"F1", x"33", x"18", x"C4", x"21", -- 0x2498,
      x"4D", x"73", x"36", x"01", x"21", x"4E", x"73", x"36", -- 0x24A0,
      x"01", x"CD", x"FE", x"17", x"21", x"61", x"28", x"E5", -- 0x24A8,
      x"21", x"C0", x"18", x"E5", x"CD", x"7C", x"06", x"F1", -- 0x24B0,
      x"F1", x"3E", x"01", x"D3", x"55", x"3E", x"0E", x"D3", -- 0x24B8,
      x"54", x"CD", x"C7", x"19", x"CD", x"8C", x"2F", x"7D", -- 0x24C0,
      x"D6", x"02", x"28", x"97", x"FD", x"21", x"48", x"73", -- 0x24C8,
      x"FD", x"7E", x"00", x"B7", x"20", x"16", x"FD", x"7E", -- 0x24D0,
      x"01", x"D6", x"80", x"20", x"0F", x"AF", x"F5", x"33", -- 0x24D8,
      x"21", x"69", x"28", x"E5", x"CD", x"F3", x"18", x"F1", -- 0x24E0,
      x"33", x"C3", x"63", x"24", x"CD", x"E3", x"1C", x"3A", -- 0x24E8,
      x"4A", x"73", x"B7", x"20", x"10", x"21", x"82", x"28", -- 0x24F0,
      x"E5", x"3E", x"01", x"F5", x"33", x"CD", x"38", x"08", -- 0x24F8,
      x"F1", x"33", x"C3", x"63", x"24", x"CD", x"FE", x"17", -- 0x2500,
      x"21", x"4B", x"73", x"36", x"00", x"21", x"4C", x"73", -- 0x2508,
      x"36", x"00", x"FD", x"21", x"4E", x"73", x"FD", x"7E", -- 0x2510,
      x"00", x"B7", x"28", x"55", x"FD", x"36", x"00", x"00", -- 0x2518,
      x"3E", x"80", x"D3", x"BF", x"3E", x"81", x"D3", x"BF", -- 0x2520,
      x"21", x"F0", x"02", x"E5", x"21", x"AF", x"14", x"E5", -- 0x2528,
      x"21", x"E8", x"08", x"E5", x"CD", x"0A", x"29", x"F1", -- 0x2530,
      x"F1", x"F1", x"FD", x"21", x"47", x"73", x"FD", x"7E", -- 0x2538,
      x"00", x"F6", x"02", x"32", x"47", x"73", x"FD", x"7E", -- 0x2540,
      x"00", x"D3", x"BF", x"3E", x"B2", x"D3", x"BF", x"3E", -- 0x2548,
      x"06", x"D3", x"BF", x"3E", x"87", x"D3", x"BF", x"CD", -- 0x2550,
      x"0F", x"18", x"21", x"38", x"72", x"36", x"00", x"CD", -- 0x2558,
      x"2B", x"24", x"3E", x"F2", x"D3", x"BF", x"3E", x"81", -- 0x2560,
      x"D3", x"BF", x"21", x"46", x"73", x"36", x"28", x"18", -- 0x2568,
      x"03", x"CD", x"0F", x"18", x"3E", x"0E", x"D3", x"54", -- 0x2570,
      x"CD", x"9D", x"1B", x"CD", x"B0", x"22", x"CB", x"7D", -- 0x2578,
      x"28", x"08", x"CD", x"9D", x"1B", x"CD", x"6C", x"1B", -- 0x2580,
      x"18", x"F1", x"CD", x"8C", x"2F", x"7D", x"D6", x"02", -- 0x2588,
      x"20", x"06", x"CD", x"0F", x"18", x"C3", x"63", x"24", -- 0x2590,
      x"FD", x"21", x"4C", x"73", x"FD", x"6E", x"00", x"26", -- 0x2598,
      x"00", x"29", x"11", x"C3", x"6A", x"19", x"4E", x"23", -- 0x25A0,
      x"46", x"69", x"60", x"11", x"7F", x"00", x"19", x"7E", -- 0x25A8,
      x"B7", x"C2", x"75", x"26", x"11", x"C3", x"66", x"1A", -- 0x25B0,
      x"B7", x"28", x"03", x"13", x"18", x"F9", x"DD", x"73", -- 0x25B8,
      x"FE", x"DD", x"72", x"FF", x"DD", x"73", x"FC", x"DD", -- 0x25C0,
      x"72", x"FD", x"0A", x"D6", x"2E", x"20", x"33", x"69", -- 0x25C8,
      x"60", x"23", x"7E", x"D6", x"2E", x"20", x"2B", x"4B", -- 0x25D0,
      x"42", x"0A", x"D6", x"2F", x"28", x"0D", x"59", x"50", -- 0x25D8,
      x"3E", x"C3", x"93", x"3E", x"66", x"9A", x"30", x"03", -- 0x25E0,
      x"0B", x"18", x"EE", x"59", x"50", x"21", x"C3", x"66", -- 0x25E8,
      x"BF", x"ED", x"52", x"20", x"09", x"36", x"2F", x"21", -- 0x25F0,
      x"C4", x"66", x"36", x"00", x"18", x"71", x"AF", x"02", -- 0x25F8,
      x"18", x"6D", x"DD", x"5E", x"FE", x"DD", x"56", x"FF", -- 0x2600,
      x"3E", x"C4", x"93", x"3E", x"66", x"9A", x"30", x"10", -- 0x2608,
      x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"36", x"2F", -- 0x2610,
      x"DD", x"34", x"FE", x"20", x"03", x"DD", x"34", x"FF", -- 0x2618,
      x"0A", x"5F", x"B7", x"28", x"29", x"DD", x"7E", x"FE", -- 0x2620,
      x"D6", x"C3", x"57", x"DD", x"7E", x"FF", x"DE", x"66", -- 0x2628,
      x"6F", x"7A", x"D6", x"FE", x"7D", x"17", x"3F", x"1F", -- 0x2630,
      x"DE", x"81", x"30", x"12", x"03", x"DD", x"6E", x"FE", -- 0x2638,
      x"DD", x"66", x"FF", x"73", x"DD", x"34", x"FE", x"20", -- 0x2640,
      x"D7", x"DD", x"34", x"FF", x"18", x"D2", x"0A", x"B7", -- 0x2648,
      x"28", x"15", x"C1", x"E1", x"E5", x"C5", x"36", x"00", -- 0x2650,
      x"AF", x"F5", x"33", x"21", x"91", x"28", x"E5", x"CD", -- 0x2658,
      x"F3", x"18", x"F1", x"33", x"C3", x"74", x"25", x"DD", -- 0x2660,
      x"6E", x"FE", x"DD", x"66", x"FF", x"36", x"00", x"CD", -- 0x2668,
      x"0F", x"18", x"C3", x"A9", x"24", x"DD", x"77", x"FD", -- 0x2670,
      x"DD", x"36", x"FE", x"C3", x"DD", x"36", x"FF", x"68", -- 0x2678,
      x"11", x"C3", x"66", x"1A", x"B7", x"28", x"12", x"13", -- 0x2680,
      x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"77", x"DD", -- 0x2688,
      x"34", x"FE", x"20", x"EF", x"DD", x"34", x"FF", x"18", -- 0x2690,
      x"EA", x"DD", x"5E", x"FE", x"DD", x"56", x"FF", x"3A", -- 0x2698,
      x"C4", x"66", x"B7", x"28", x"0F", x"DD", x"6E", x"FE", -- 0x26A0,
      x"DD", x"66", x"FF", x"36", x"2F", x"DD", x"5E", x"FE", -- 0x26A8,
      x"DD", x"56", x"FF", x"13", x"0A", x"DD", x"77", x"FF", -- 0x26B0,
      x"B7", x"28", x"1B", x"7B", x"D6", x"C3", x"6F", x"7A", -- 0x26B8,
      x"DE", x"68", x"67", x"7D", x"D6", x"7F", x"7C", x"17", -- 0x26C0,
      x"3F", x"1F", x"DE", x"80", x"30", x"08", x"DD", x"7E", -- 0x26C8,
      x"FF", x"03", x"12", x"13", x"18", x"DE", x"AF", x"12", -- 0x26D0,
      x"0A", x"B7", x"28", x"10", x"3E", x"01", x"F5", x"33", -- 0x26D8,
      x"21", x"91", x"28", x"E5", x"CD", x"F3", x"18", x"F1", -- 0x26E0,
      x"33", x"C3", x"74", x"25", x"CD", x"22", x"18", x"21", -- 0x26E8,
      x"A2", x"28", x"E5", x"AF", x"F5", x"33", x"CD", x"38", -- 0x26F0,
      x"08", x"33", x"21", x"C3", x"68", x"E3", x"21", x"EC", -- 0x26F8,
      x"6E", x"E5", x"CD", x"8D", x"30", x"F1", x"F1", x"45", -- 0x2700,
      x"78", x"B7", x"28", x"0E", x"C5", x"33", x"21", x"AE", -- 0x2708,
      x"28", x"E5", x"CD", x"F3", x"18", x"F1", x"33", x"C3", -- 0x2710,
      x"74", x"25", x"3E", x"01", x"D3", x"54", x"21", x"00", -- 0x2718,
      x"00", x"39", x"4D", x"44", x"59", x"50", x"C5", x"D5", -- 0x2720,
      x"21", x"00", x"02", x"E5", x"26", x"80", x"E5", x"21", -- 0x2728,
      x"EC", x"6E", x"E5", x"CD", x"DC", x"29", x"F1", x"F1", -- 0x2730,
      x"F1", x"F1", x"C1", x"DD", x"75", x"FF", x"7D", x"B7", -- 0x2738,
      x"20", x"0D", x"DD", x"7E", x"FA", x"B7", x"20", x"07", -- 0x2740,
      x"DD", x"7E", x"FB", x"D6", x"02", x"28", x"19", x"21", -- 0x2748,
      x"EC", x"6E", x"E5", x"CD", x"7B", x"46", x"F1", x"DD", -- 0x2750,
      x"7E", x"FF", x"F5", x"33", x"21", x"C3", x"28", x"E5", -- 0x2758,
      x"CD", x"F3", x"18", x"F1", x"33", x"C3", x"74", x"25", -- 0x2760,
      x"3A", x"00", x"80", x"D6", x"AA", x"20", x"07", x"3A", -- 0x2768,
      x"01", x"80", x"D6", x"55", x"28", x"0E", x"3A", x"00", -- 0x2770,
      x"80", x"D6", x"55", x"20", x"0D", x"3A", x"01", x"80", -- 0x2778,
      x"D6", x"AA", x"20", x"06", x"CD", x"AF", x"1E", x"C3", -- 0x2780,
      x"74", x"25", x"DD", x"6E", x"FD", x"26", x"00", x"2B", -- 0x2788,
      x"7C", x"17", x"9F", x"5F", x"57", x"3E", x"0E", x"29", -- 0x2790,
      x"CB", x"13", x"CB", x"12", x"3D", x"20", x"F8", x"C5", -- 0x2798,
      x"D5", x"E5", x"21", x"EC", x"6E", x"E5", x"CD", x"46", -- 0x27A0,
      x"3F", x"F1", x"F1", x"F1", x"7D", x"C1", x"B7", x"28", -- 0x27A8,
      x"19", x"21", x"EC", x"6E", x"E5", x"CD", x"7B", x"46", -- 0x27B0,
      x"F1", x"DD", x"7E", x"FF", x"F5", x"33", x"21", x"DB", -- 0x27B8,
      x"28", x"E5", x"CD", x"F3", x"18", x"F1", x"33", x"C3", -- 0x27C0,
      x"74", x"25", x"C5", x"21", x"00", x"02", x"E5", x"26", -- 0x27C8,
      x"82", x"E5", x"21", x"EC", x"6E", x"E5", x"CD", x"DC", -- 0x27D0,
      x"29", x"F1", x"F1", x"F1", x"F1", x"4D", x"79", x"B7", -- 0x27D8,
      x"20", x"0D", x"DD", x"7E", x"FA", x"B7", x"20", x"07", -- 0x27E0,
      x"DD", x"7E", x"FB", x"D6", x"02", x"28", x"19", x"C5", -- 0x27E8,
      x"21", x"EC", x"6E", x"E5", x"CD", x"7B", x"46", x"F1", -- 0x27F0,
      x"C1", x"79", x"F5", x"33", x"21", x"F4", x"28", x"E5", -- 0x27F8,
      x"CD", x"F3", x"18", x"F1", x"33", x"C3", x"74", x"25", -- 0x2800,
      x"3A", x"00", x"82", x"D6", x"AA", x"20", x"07", x"3A", -- 0x2808,
      x"01", x"82", x"D6", x"55", x"28", x"0E", x"3A", x"00", -- 0x2810,
      x"82", x"D6", x"55", x"20", x"19", x"3A", x"01", x"82", -- 0x2818,
      x"D6", x"AA", x"20", x"12", x"DD", x"7E", x"FD", x"F5", -- 0x2820,
      x"33", x"CD", x"E1", x"1F", x"33", x"7D", x"D6", x"0E", -- 0x2828,
      x"DA", x"74", x"25", x"C3", x"A9", x"24", x"21", x"EC", -- 0x2830,
      x"6E", x"E5", x"CD", x"7B", x"46", x"F1", x"AF", x"F5", -- 0x2838,
      x"33", x"21", x"C3", x"28", x"E5", x"CD", x"F3", x"18", -- 0x2840,
      x"F1", x"33", x"C3", x"74", x"25", x"00", x"46", x"61", -- 0x2848,
      x"69", x"6C", x"65", x"64", x"20", x"74", x"6F", x"20", -- 0x2850,
      x"6D", x"6F", x"75", x"6E", x"74", x"20", x"53", x"44", -- 0x2858,
      x"00", x"52", x"45", x"41", x"44", x"49", x"4E", x"47", -- 0x2860,
      x"00", x"46", x"61", x"69", x"6C", x"65", x"64", x"20", -- 0x2868,
      x"74", x"6F", x"20", x"6F", x"70", x"65", x"6E", x"20", -- 0x2870,
      x"64", x"69", x"72", x"65", x"63", x"74", x"6F", x"72", -- 0x2878,
      x"79", x"00", x"4E", x"6F", x"20", x"66", x"69", x"6C", -- 0x2880,
      x"65", x"73", x"20", x"66", x"6F", x"75", x"6E", x"64", -- 0x2888,
      x"00", x"50", x"61", x"74", x"68", x"20", x"74", x"6F", -- 0x2890,
      x"6F", x"20", x"6C", x"6F", x"6E", x"67", x"2E", x"2E", -- 0x2898,
      x"2E", x"00", x"63", x"68", x"65", x"63", x"6B", x"69", -- 0x28A0,
      x"6E", x"67", x"2E", x"2E", x"2E", x"00", x"46", x"61", -- 0x28A8,
      x"69", x"6C", x"65", x"64", x"20", x"74", x"6F", x"20", -- 0x28B0,
      x"6F", x"70", x"65", x"6E", x"20", x"66", x"69", x"6C", -- 0x28B8,
      x"65", x"2E", x"00", x"55", x"6E", x"72", x"65", x"63", -- 0x28C0,
      x"6F", x"67", x"6E", x"69", x"7A", x"65", x"64", x"20", -- 0x28C8,
      x"66", x"69", x"6C", x"65", x"20", x"74", x"79", x"70", -- 0x28D0,
      x"65", x"2E", x"00", x"46", x"61", x"69", x"6C", x"65", -- 0x28D8,
      x"64", x"20", x"74", x"6F", x"20", x"69", x"64", x"65", -- 0x28E0,
      x"6E", x"74", x"69", x"66", x"79", x"20", x"66", x"69", -- 0x28E8,
      x"6C", x"65", x"2E", x"00", x"46", x"61", x"69", x"6C", -- 0x28F0,
      x"65", x"64", x"20", x"74", x"6F", x"20", x"72", x"65", -- 0x28F8,
      x"61", x"64", x"20", x"62", x"6C", x"6F", x"63", x"6B", -- 0x2900,
      x"2E", x"00", x"DD", x"E5", x"E5", x"C5", x"D5", x"F5", -- 0x2908,
      x"DD", x"21", x"0C", x"00", x"DD", x"39", x"DD", x"5E", -- 0x2910,
      x"00", x"DD", x"56", x"01", x"7B", x"D3", x"BF", x"7A", -- 0x2918,
      x"CB", x"F7", x"D3", x"BF", x"DD", x"6E", x"02", x"DD", -- 0x2920,
      x"66", x"03", x"DD", x"5E", x"04", x"DD", x"56", x"05", -- 0x2928,
      x"0E", x"BE", x"14", x"15", x"28", x"07", x"AF", x"47", -- 0x2930,
      x"ED", x"B3", x"15", x"18", x"F5", x"1C", x"1D", x"28", -- 0x2938,
      x"03", x"43", x"ED", x"B3", x"F1", x"D1", x"C1", x"E1", -- 0x2940,
      x"DD", x"E1", x"C9", x"CD", x"13", x"3F", x"3E", x"2A", -- 0x2948,
      x"D3", x"80", x"DD", x"7E", x"04", x"D6", x"02", x"3E", -- 0x2950,
      x"01", x"28", x"01", x"AF", x"4F", x"B7", x"28", x"05", -- 0x2958,
      x"DB", x"FF", x"5F", x"18", x"03", x"DB", x"FC", x"5F", -- 0x2960,
      x"CB", x"73", x"20", x"07", x"21", x"39", x"72", x"36", -- 0x2968,
      x"12", x"18", x"0F", x"7B", x"E6", x"0F", x"5F", x"16", -- 0x2970,
      x"00", x"21", x"CC", x"29", x"19", x"EB", x"1A", x"32", -- 0x2978,
      x"39", x"72", x"21", x"3B", x"72", x"36", x"00", x"21", -- 0x2980,
      x"3A", x"72", x"36", x"00", x"3E", x"2A", x"D3", x"C0", -- 0x2988,
      x"79", x"B7", x"28", x"05", x"DB", x"FF", x"4F", x"18", -- 0x2990,
      x"03", x"DB", x"FC", x"4F", x"CB", x"71", x"20", x"05", -- 0x2998,
      x"21", x"39", x"72", x"36", x"12", x"CB", x"59", x"20", -- 0x29A0,
      x"05", x"21", x"3B", x"72", x"36", x"FC", x"CB", x"51", -- 0x29A8,
      x"20", x"05", x"21", x"3A", x"72", x"36", x"FC", x"CB", -- 0x29B0,
      x"49", x"20", x"05", x"21", x"3B", x"72", x"36", x"04", -- 0x29B8,
      x"CB", x"41", x"20", x"05", x"21", x"3A", x"72", x"36", -- 0x29C0,
      x"04", x"DD", x"E1", x"C9", x"FF", x"38", x"34", x"35", -- 0x29C8,
      x"FF", x"37", x"23", x"32", x"FF", x"2A", x"30", x"39", -- 0x29D0,
      x"33", x"31", x"36", x"FF", x"CD", x"13", x"3F", x"21", -- 0x29D8,
      x"E0", x"FF", x"39", x"F9", x"DD", x"7E", x"06", x"DD", -- 0x29E0,
      x"77", x"FE", x"DD", x"7E", x"07", x"DD", x"77", x"FF", -- 0x29E8,
      x"DD", x"7E", x"0A", x"DD", x"77", x"E2", x"DD", x"7E", -- 0x29F0,
      x"0B", x"DD", x"77", x"E3", x"C1", x"E1", x"E5", x"C5", -- 0x29F8,
      x"AF", x"77", x"23", x"77", x"21", x"00", x"00", x"39", -- 0x2A00,
      x"DD", x"7E", x"04", x"DD", x"77", x"E4", x"DD", x"7E", -- 0x2A08,
      x"05", x"DD", x"77", x"E5", x"E5", x"DD", x"6E", x"E4", -- 0x2A10,
      x"DD", x"66", x"E5", x"E5", x"CD", x"A5", x"35", x"F1", -- 0x2A18,
      x"F1", x"4D", x"DD", x"71", x"FD", x"79", x"B7", x"20", -- 0x2A20,
      x"1D", x"DD", x"7E", x"E4", x"C6", x"0F", x"DD", x"77", -- 0x2A28,
      x"E6", x"DD", x"7E", x"E5", x"CE", x"00", x"DD", x"77", -- 0x2A30,
      x"E7", x"DD", x"6E", x"E6", x"DD", x"66", x"E7", x"7E", -- 0x2A38,
      x"DD", x"77", x"FD", x"B7", x"28", x"06", x"DD", x"6E", -- 0x2A40,
      x"FD", x"C3", x"26", x"2E", x"DD", x"7E", x"E4", x"DD", -- 0x2A48,
      x"77", x"E8", x"DD", x"7E", x"E5", x"DD", x"77", x"E9", -- 0x2A50,
      x"DD", x"6E", x"E4", x"DD", x"66", x"E5", x"11", x"0E", -- 0x2A58,
      x"00", x"19", x"7E", x"0F", x"38", x"05", x"2E", x"07", -- 0x2A60,
      x"C3", x"26", x"2E", x"DD", x"6E", x"E4", x"DD", x"66", -- 0x2A68,
      x"E5", x"11", x"0A", x"00", x"19", x"4E", x"23", x"46", -- 0x2A70,
      x"23", x"5E", x"23", x"56", x"DD", x"7E", x"E4", x"C6", -- 0x2A78,
      x"10", x"DD", x"77", x"EA", x"DD", x"7E", x"E5", x"CE", -- 0x2A80,
      x"00", x"DD", x"77", x"EB", x"D5", x"C5", x"DD", x"5E", -- 0x2A88,
      x"EA", x"DD", x"56", x"EB", x"21", x"1E", x"00", x"39", -- 0x2A90,
      x"EB", x"01", x"04", x"00", x"ED", x"B0", x"C1", x"D1", -- 0x2A98,
      x"79", x"DD", x"96", x"FA", x"4F", x"78", x"DD", x"9E", -- 0x2AA0,
      x"FB", x"47", x"7B", x"DD", x"9E", x"FC", x"5F", x"7A", -- 0x2AA8,
      x"DD", x"9E", x"FD", x"57", x"DD", x"7E", x"08", x"DD", -- 0x2AB0,
      x"77", x"FA", x"DD", x"7E", x"09", x"DD", x"77", x"FB", -- 0x2AB8,
      x"AF", x"DD", x"77", x"FC", x"DD", x"77", x"FD", x"79", -- 0x2AC0,
      x"DD", x"96", x"FA", x"78", x"DD", x"9E", x"FB", x"7B", -- 0x2AC8,
      x"DD", x"9E", x"FC", x"7A", x"DD", x"9E", x"FD", x"30", -- 0x2AD0,
      x"06", x"DD", x"71", x"08", x"DD", x"70", x"09", x"DD", -- 0x2AD8,
      x"7E", x"E4", x"DD", x"77", x"EC", x"DD", x"7E", x"E5", -- 0x2AE0,
      x"DD", x"77", x"ED", x"DD", x"7E", x"E4", x"DD", x"77", -- 0x2AE8,
      x"EE", x"DD", x"7E", x"E5", x"DD", x"77", x"EF", x"DD", -- 0x2AF0,
      x"7E", x"EA", x"DD", x"77", x"F0", x"DD", x"7E", x"EB", -- 0x2AF8,
      x"DD", x"77", x"F1", x"DD", x"7E", x"E4", x"C6", x"1C", -- 0x2B00,
      x"DD", x"77", x"F2", x"DD", x"7E", x"E5", x"CE", x"00", -- 0x2B08,
      x"DD", x"77", x"F3", x"DD", x"7E", x"E4", x"DD", x"77", -- 0x2B10,
      x"F4", x"DD", x"7E", x"E5", x"DD", x"77", x"F5", x"DD", -- 0x2B18,
      x"7E", x"09", x"DD", x"B6", x"08", x"CA", x"24", x"2E", -- 0x2B20,
      x"DD", x"6E", x"EA", x"DD", x"66", x"EB", x"4E", x"23", -- 0x2B28,
      x"46", x"23", x"5E", x"23", x"56", x"79", x"B7", x"C2", -- 0x2B30,
      x"5A", x"2D", x"CB", x"40", x"C2", x"5A", x"2D", x"DD", -- 0x2B38,
      x"70", x"FA", x"DD", x"73", x"FB", x"DD", x"72", x"FC", -- 0x2B40,
      x"AF", x"DD", x"77", x"FD", x"DD", x"CB", x"FC", x"3E", -- 0x2B48,
      x"DD", x"CB", x"FB", x"1E", x"DD", x"CB", x"FA", x"1E", -- 0x2B50,
      x"E1", x"E5", x"C5", x"01", x"09", x"00", x"09", x"C1", -- 0x2B58,
      x"7E", x"2B", x"6E", x"67", x"2B", x"DD", x"7E", x"FA", -- 0x2B60,
      x"DD", x"77", x"FC", x"DD", x"7E", x"FB", x"DD", x"77", -- 0x2B68,
      x"FD", x"7D", x"DD", x"A6", x"FC", x"6F", x"7C", x"DD", -- 0x2B70,
      x"A6", x"FD", x"67", x"DD", x"75", x"FC", x"DD", x"74", -- 0x2B78,
      x"FD", x"7C", x"DD", x"B6", x"FC", x"C2", x"11", x"2C", -- 0x2B80,
      x"7A", x"B3", x"B0", x"B1", x"20", x"13", x"DD", x"6E", -- 0x2B88,
      x"EC", x"DD", x"66", x"ED", x"11", x"06", x"00", x"19", -- 0x2B90,
      x"4E", x"23", x"46", x"23", x"5E", x"23", x"56", x"18", -- 0x2B98,
      x"2E", x"DD", x"7E", x"E8", x"DD", x"77", x"FA", x"DD", -- 0x2BA0,
      x"7E", x"E9", x"DD", x"77", x"FB", x"DD", x"6E", x"FA", -- 0x2BA8,
      x"DD", x"66", x"FB", x"11", x"14", x"00", x"19", x"4E", -- 0x2BB0,
      x"23", x"46", x"23", x"5E", x"23", x"56", x"D5", x"C5", -- 0x2BB8,
      x"DD", x"6E", x"E8", x"DD", x"66", x"E9", x"E5", x"CD", -- 0x2BC0,
      x"C1", x"44", x"F1", x"F1", x"F1", x"4D", x"44", x"79", -- 0x2BC8,
      x"D6", x"02", x"78", x"DE", x"00", x"7B", x"DE", x"00", -- 0x2BD0,
      x"7A", x"DE", x"00", x"30", x"0D", x"DD", x"6E", x"E6", -- 0x2BD8,
      x"DD", x"66", x"E7", x"36", x"02", x"2E", x"02", x"C3", -- 0x2BE0,
      x"26", x"2E", x"79", x"A0", x"A3", x"A2", x"3C", x"20", -- 0x2BE8,
      x"0D", x"DD", x"6E", x"E6", x"DD", x"66", x"E7", x"36", -- 0x2BF0,
      x"01", x"2E", x"01", x"C3", x"26", x"2E", x"DD", x"7E", -- 0x2BF8,
      x"EE", x"C6", x"14", x"6F", x"DD", x"7E", x"EF", x"CE", -- 0x2C00,
      x"00", x"67", x"71", x"23", x"70", x"23", x"73", x"23", -- 0x2C08,
      x"72", x"DD", x"6E", x"E4", x"DD", x"66", x"E5", x"11", -- 0x2C10,
      x"14", x"00", x"19", x"4E", x"23", x"46", x"23", x"5E", -- 0x2C18,
      x"23", x"56", x"D5", x"C5", x"DD", x"6E", x"E0", x"DD", -- 0x2C20,
      x"66", x"E1", x"E5", x"CD", x"68", x"37", x"F1", x"F1", -- 0x2C28,
      x"F1", x"7A", x"B3", x"B4", x"B5", x"20", x"0D", x"DD", -- 0x2C30,
      x"6E", x"E6", x"DD", x"66", x"E7", x"36", x"02", x"2E", -- 0x2C38,
      x"02", x"C3", x"26", x"2E", x"DD", x"7E", x"FC", x"DD", -- 0x2C40,
      x"77", x"F8", x"DD", x"7E", x"FD", x"DD", x"77", x"F9", -- 0x2C48,
      x"AF", x"DD", x"77", x"FA", x"DD", x"77", x"FB", x"7D", -- 0x2C50,
      x"DD", x"86", x"F8", x"4F", x"7C", x"DD", x"8E", x"F9", -- 0x2C58,
      x"47", x"7B", x"DD", x"8E", x"FA", x"5F", x"7A", x"DD", -- 0x2C60,
      x"8E", x"FB", x"57", x"DD", x"71", x"F8", x"DD", x"70", -- 0x2C68,
      x"F9", x"DD", x"73", x"FA", x"DD", x"72", x"FB", x"DD", -- 0x2C70,
      x"7E", x"09", x"CB", x"3F", x"4F", x"06", x"00", x"78", -- 0x2C78,
      x"B1", x"28", x"5D", x"DD", x"7E", x"FC", x"81", x"5F", -- 0x2C80,
      x"DD", x"7E", x"FD", x"88", x"57", x"E1", x"E5", x"C5", -- 0x2C88,
      x"01", x"08", x"00", x"09", x"C1", x"7E", x"23", x"66", -- 0x2C90,
      x"6F", x"93", x"7C", x"9A", x"30", x"0A", x"7D", x"DD", -- 0x2C98,
      x"96", x"FC", x"4F", x"7C", x"DD", x"9E", x"FD", x"47", -- 0x2CA0,
      x"C5", x"C5", x"DD", x"6E", x"FA", x"DD", x"66", x"FB", -- 0x2CA8,
      x"E5", x"DD", x"6E", x"F8", x"DD", x"66", x"F9", x"E5", -- 0x2CB0,
      x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"E5", x"CD", -- 0x2CB8,
      x"61", x"2E", x"F1", x"F1", x"F1", x"F1", x"7D", x"C1", -- 0x2CC0,
      x"B7", x"28", x"0D", x"DD", x"6E", x"E6", x"DD", x"66", -- 0x2CC8,
      x"E7", x"36", x"01", x"2E", x"01", x"C3", x"26", x"2E", -- 0x2CD0,
      x"79", x"87", x"47", x"0E", x"00", x"C3", x"AE", x"2D", -- 0x2CD8,
      x"DD", x"7E", x"E4", x"C6", x"18", x"DD", x"77", x"FC", -- 0x2CE0,
      x"DD", x"7E", x"E5", x"CE", x"00", x"DD", x"77", x"FD", -- 0x2CE8,
      x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"4E", x"23", -- 0x2CF0,
      x"46", x"23", x"5E", x"23", x"56", x"DD", x"7E", x"F8", -- 0x2CF8,
      x"91", x"20", x"11", x"DD", x"7E", x"F9", x"90", x"20", -- 0x2D00,
      x"0B", x"DD", x"6E", x"FA", x"DD", x"66", x"FB", x"BF", -- 0x2D08,
      x"ED", x"52", x"28", x"37", x"DD", x"7E", x"E4", x"C6", -- 0x2D10,
      x"1C", x"4F", x"DD", x"7E", x"E5", x"CE", x"00", x"47", -- 0x2D18,
      x"21", x"01", x"00", x"E5", x"DD", x"6E", x"FA", x"DD", -- 0x2D20,
      x"66", x"FB", x"E5", x"DD", x"6E", x"F8", x"DD", x"66", -- 0x2D28,
      x"F9", x"E5", x"C5", x"CD", x"61", x"2E", x"F1", x"F1", -- 0x2D30,
      x"F1", x"F1", x"7D", x"B7", x"28", x"0D", x"DD", x"6E", -- 0x2D38,
      x"E6", x"DD", x"66", x"E7", x"36", x"01", x"2E", x"01", -- 0x2D40,
      x"C3", x"26", x"2E", x"DD", x"5E", x"FC", x"DD", x"56", -- 0x2D48,
      x"FD", x"21", x"18", x"00", x"39", x"01", x"04", x"00", -- 0x2D50,
      x"ED", x"B0", x"DD", x"5E", x"F0", x"DD", x"56", x"F1", -- 0x2D58,
      x"21", x"1A", x"00", x"39", x"EB", x"01", x"04", x"00", -- 0x2D60,
      x"ED", x"B0", x"DD", x"4E", x"FA", x"DD", x"7E", x"FB", -- 0x2D68,
      x"E6", x"01", x"47", x"AF", x"91", x"4F", x"3E", x"02", -- 0x2D70,
      x"98", x"47", x"DD", x"7E", x"08", x"91", x"DD", x"7E", -- 0x2D78,
      x"09", x"98", x"30", x"06", x"DD", x"4E", x"08", x"DD", -- 0x2D80,
      x"46", x"09", x"DD", x"5E", x"FA", x"DD", x"7E", x"FB", -- 0x2D88,
      x"E6", x"01", x"57", x"7B", x"DD", x"86", x"F2", x"5F", -- 0x2D90,
      x"7A", x"DD", x"8E", x"F3", x"57", x"DD", x"6E", x"FE", -- 0x2D98,
      x"DD", x"66", x"FF", x"C5", x"C5", x"D5", x"E5", x"CD", -- 0x2DA0,
      x"AE", x"00", x"F1", x"F1", x"F1", x"C1", x"DD", x"7E", -- 0x2DA8,
      x"08", x"91", x"DD", x"77", x"08", x"DD", x"7E", x"09", -- 0x2DB0,
      x"98", x"DD", x"77", x"09", x"DD", x"6E", x"E2", x"DD", -- 0x2DB8,
      x"66", x"E3", x"7E", x"23", x"66", x"6F", x"09", x"EB", -- 0x2DC0,
      x"DD", x"6E", x"E2", x"DD", x"66", x"E3", x"73", x"23", -- 0x2DC8,
      x"72", x"DD", x"7E", x"FE", x"81", x"DD", x"77", x"FE", -- 0x2DD0,
      x"DD", x"7E", x"FF", x"88", x"DD", x"77", x"FF", x"DD", -- 0x2DD8,
      x"7E", x"F4", x"C6", x"10", x"5F", x"DD", x"7E", x"F5", -- 0x2DE0,
      x"CE", x"00", x"57", x"D5", x"C5", x"21", x"1A", x"00", -- 0x2DE8,
      x"39", x"EB", x"01", x"04", x"00", x"ED", x"B0", x"C1", -- 0x2DF0,
      x"D1", x"21", x"00", x"00", x"79", x"DD", x"86", x"F6", -- 0x2DF8,
      x"DD", x"77", x"FA", x"78", x"DD", x"8E", x"F7", x"DD", -- 0x2E00,
      x"77", x"FB", x"7D", x"DD", x"8E", x"F8", x"DD", x"77", -- 0x2E08,
      x"FC", x"7C", x"DD", x"8E", x"F9", x"DD", x"77", x"FD", -- 0x2E10,
      x"21", x"1A", x"00", x"39", x"01", x"04", x"00", x"ED", -- 0x2E18,
      x"B0", x"C3", x"1F", x"2B", x"2E", x"00", x"DD", x"F9", -- 0x2E20,
      x"DD", x"E1", x"C9", x"DD", x"E5", x"DD", x"21", x"00", -- 0x2E28,
      x"00", x"DD", x"39", x"DD", x"7E", x"04", x"DD", x"4E", -- 0x2E30,
      x"05", x"D3", x"BF", x"06", x"00", x"79", x"D3", x"BF", -- 0x2E38,
      x"00", x"00", x"00", x"00", x"00", x"DD", x"4E", x"06", -- 0x2E40,
      x"DD", x"46", x"07", x"DD", x"5E", x"08", x"DD", x"56", -- 0x2E48,
      x"09", x"6B", x"62", x"1B", x"7C", x"B5", x"28", x"06", -- 0x2E50,
      x"DB", x"BE", x"02", x"03", x"18", x"F3", x"DD", x"E1", -- 0x2E58,
      x"C9", x"CD", x"13", x"3F", x"F5", x"3B", x"CD", x"8C", -- 0x2E60,
      x"2F", x"7D", x"0F", x"30", x"05", x"2E", x"03", x"C3", -- 0x2E68,
      x"22", x"2F", x"3A", x"3E", x"72", x"CB", x"5F", x"20", -- 0x2E70,
      x"14", x"06", x"09", x"DD", x"CB", x"06", x"26", x"DD", -- 0x2E78,
      x"CB", x"07", x"16", x"DD", x"CB", x"08", x"16", x"DD", -- 0x2E80,
      x"CB", x"09", x"16", x"10", x"EE", x"3E", x"01", x"DD", -- 0x2E88,
      x"BE", x"0A", x"3E", x"00", x"DD", x"9E", x"0B", x"30", -- 0x2E90,
      x"04", x"3E", x"12", x"18", x"02", x"3E", x"11", x"DD", -- 0x2E98,
      x"77", x"FD", x"DD", x"6E", x"08", x"DD", x"66", x"09", -- 0x2EA0,
      x"E5", x"DD", x"6E", x"06", x"DD", x"66", x"07", x"E5", -- 0x2EA8,
      x"DD", x"7E", x"FD", x"F5", x"33", x"CD", x"31", x"32", -- 0x2EB0,
      x"F1", x"F1", x"33", x"7D", x"B7", x"20", x"50", x"DD", -- 0x2EB8,
      x"6E", x"04", x"DD", x"66", x"05", x"DD", x"4E", x"0A", -- 0x2EC0,
      x"DD", x"46", x"0B", x"E5", x"C5", x"11", x"00", x"02", -- 0x2EC8,
      x"D5", x"E5", x"CD", x"76", x"33", x"F1", x"F1", x"DD", -- 0x2ED0,
      x"75", x"FE", x"DD", x"74", x"FF", x"C1", x"E1", x"DD", -- 0x2ED8,
      x"7E", x"FF", x"DD", x"B6", x"FE", x"28", x"09", x"11", -- 0x2EE0,
      x"00", x"02", x"19", x"0B", x"78", x"B1", x"20", x"DB", -- 0x2EE8,
      x"DD", x"71", x"0A", x"DD", x"70", x"0B", x"DD", x"7E", -- 0x2EF0,
      x"FD", x"D6", x"12", x"20", x"12", x"21", x"00", x"00", -- 0x2EF8,
      x"E5", x"21", x"00", x"00", x"E5", x"3E", x"0C", x"F5", -- 0x2F00,
      x"33", x"CD", x"31", x"32", x"F1", x"F1", x"33", x"CD", -- 0x2F08,
      x"8F", x"35", x"DD", x"7E", x"0B", x"DD", x"B6", x"0A", -- 0x2F10,
      x"28", x"05", x"21", x"01", x"00", x"18", x"03", x"21", -- 0x2F18,
      x"00", x"00", x"DD", x"F9", x"DD", x"E1", x"C9", x"21", -- 0x2F20,
      x"43", x"73", x"36", x"00", x"DB", x"BF", x"32", x"56", -- 0x2F28,
      x"73", x"3A", x"59", x"73", x"3C", x"32", x"59", x"73", -- 0x2F30,
      x"FD", x"21", x"57", x"73", x"FD", x"7E", x"01", x"FD", -- 0x2F38,
      x"B6", x"00", x"C8", x"2A", x"57", x"73", x"E9", x"FD", -- 0x2F40,
      x"21", x"02", x"00", x"FD", x"39", x"FD", x"7E", x"00", -- 0x2F48,
      x"32", x"57", x"73", x"FD", x"7E", x"01", x"32", x"58", -- 0x2F50,
      x"73", x"C9", x"21", x"00", x"00", x"22", x"57", x"73", -- 0x2F58,
      x"C9", x"F5", x"3E", x"9F", x"D3", x"FF", x"3E", x"BF", -- 0x2F60,
      x"D3", x"FF", x"3E", x"DF", x"D3", x"FF", x"3E", x"FF", -- 0x2F68,
      x"D3", x"FF", x"21", x"43", x"73", x"36", x"00", x"21", -- 0x2F70,
      x"60", x"EA", x"E3", x"C1", x"C5", x"03", x"33", x"33", -- 0x2F78,
      x"C5", x"78", x"B1", x"20", x"F6", x"DB", x"BF", x"32", -- 0x2F80,
      x"56", x"73", x"F1", x"C9", x"DB", x"56", x"07", x"30", -- 0x2F88,
      x"08", x"FD", x"21", x"5A", x"73", x"FD", x"6E", x"00", -- 0x2F90,
      x"C9", x"2E", x"02", x"C9", x"CD", x"13", x"3F", x"F5", -- 0x2F98,
      x"F5", x"F5", x"F5", x"DD", x"7E", x"05", x"DD", x"B6", -- 0x2FA0,
      x"04", x"20", x"05", x"2E", x"09", x"C3", x"88", x"30", -- 0x2FA8,
      x"21", x"00", x"00", x"39", x"E5", x"CD", x"20", x"38", -- 0x2FB0,
      x"F1", x"4D", x"DD", x"5E", x"04", x"DD", x"56", x"05", -- 0x2FB8,
      x"79", x"B7", x"C2", x"7F", x"30", x"6B", x"62", x"DD", -- 0x2FC0,
      x"7E", x"F8", x"77", x"23", x"DD", x"7E", x"F9", x"77", -- 0x2FC8,
      x"D5", x"DD", x"6E", x"06", x"DD", x"66", x"07", x"E5", -- 0x2FD0,
      x"D5", x"CD", x"CA", x"49", x"F1", x"F1", x"7D", x"D1", -- 0x2FD8,
      x"4F", x"B7", x"C2", x"78", x"30", x"6B", x"62", x"C5", -- 0x2FE0,
      x"01", x"27", x"00", x"09", x"C1", x"7E", x"07", x"38", -- 0x2FE8,
      x"54", x"6B", x"62", x"23", x"23", x"23", x"23", x"CB", -- 0x2FF0,
      x"66", x"28", x"48", x"21", x"06", x"00", x"19", x"DD", -- 0x2FF8,
      x"75", x"FA", x"DD", x"74", x"FB", x"6B", x"62", x"C5", -- 0x3000,
      x"01", x"1A", x"00", x"09", x"C1", x"46", x"23", x"66", -- 0x3008,
      x"C5", x"D5", x"68", x"E5", x"DD", x"6E", x"F8", x"DD", -- 0x3010,
      x"66", x"F9", x"E5", x"CD", x"38", x"44", x"F1", x"F1", -- 0x3018,
      x"DD", x"75", x"FC", x"DD", x"74", x"FD", x"DD", x"73", -- 0x3020,
      x"FE", x"DD", x"72", x"FF", x"D1", x"C1", x"D5", x"C5", -- 0x3028,
      x"DD", x"5E", x"FA", x"DD", x"56", x"FB", x"21", x"08", -- 0x3030,
      x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", x"C1", -- 0x3038,
      x"D1", x"18", x"02", x"0E", x"05", x"79", x"B7", x"20", -- 0x3040,
      x"2F", x"21", x"02", x"00", x"19", x"DD", x"75", x"FE", -- 0x3048,
      x"DD", x"74", x"FF", x"E1", x"E5", x"01", x"04", x"00", -- 0x3050,
      x"09", x"4E", x"23", x"46", x"DD", x"6E", x"FE", x"DD", -- 0x3058,
      x"66", x"FF", x"71", x"23", x"70", x"D5", x"21", x"00", -- 0x3060,
      x"00", x"E5", x"21", x"00", x"00", x"E5", x"D5", x"CD", -- 0x3068,
      x"B6", x"46", x"F1", x"F1", x"F1", x"7D", x"D1", x"4F", -- 0x3070,
      x"79", x"D6", x"04", x"20", x"02", x"0E", x"05", x"79", -- 0x3078,
      x"B7", x"28", x"04", x"AF", x"12", x"13", x"12", x"69", -- 0x3080,
      x"DD", x"F9", x"DD", x"E1", x"C9", x"CD", x"13", x"3F", -- 0x3088,
      x"21", x"CB", x"FF", x"39", x"F9", x"DD", x"7E", x"05", -- 0x3090,
      x"DD", x"B6", x"04", x"20", x"05", x"2E", x"09", x"C3", -- 0x3098,
      x"ED", x"31", x"21", x"2C", x"00", x"39", x"E5", x"CD", -- 0x30A0,
      x"20", x"38", x"F1", x"DD", x"75", x"F9", x"DD", x"4E", -- 0x30A8,
      x"04", x"DD", x"46", x"05", x"DD", x"7E", x"F9", x"B7", -- 0x30B0,
      x"C2", x"E0", x"31", x"21", x"00", x"00", x"39", x"DD", -- 0x30B8,
      x"7E", x"F7", x"77", x"23", x"DD", x"7E", x"F8", x"77", -- 0x30C0,
      x"21", x"00", x"00", x"39", x"EB", x"DD", x"73", x"FE", -- 0x30C8,
      x"DD", x"72", x"FF", x"C5", x"D5", x"DD", x"6E", x"06", -- 0x30D0,
      x"DD", x"66", x"07", x"E5", x"DD", x"6E", x"FE", x"DD", -- 0x30D8,
      x"66", x"FF", x"E5", x"CD", x"CA", x"49", x"F1", x"F1", -- 0x30E0,
      x"D1", x"C1", x"DD", x"75", x"F9", x"7D", x"B7", x"20", -- 0x30E8,
      x"20", x"6B", x"62", x"C5", x"01", x"27", x"00", x"09", -- 0x30F0,
      x"C1", x"7E", x"07", x"30", x"06", x"DD", x"36", x"F9", -- 0x30F8,
      x"06", x"18", x"0E", x"6B", x"62", x"23", x"23", x"23", -- 0x3100,
      x"23", x"CB", x"66", x"28", x"04", x"DD", x"36", x"F9", -- 0x3108,
      x"04", x"DD", x"7E", x"F9", x"B7", x"C2", x"E0", x"31", -- 0x3110,
      x"21", x"06", x"00", x"09", x"DD", x"75", x"FA", x"DD", -- 0x3118,
      x"74", x"FB", x"21", x"1A", x"00", x"19", x"EB", x"6B", -- 0x3120,
      x"62", x"7E", x"23", x"66", x"6F", x"C5", x"D5", x"E5", -- 0x3128,
      x"DD", x"6E", x"F7", x"DD", x"66", x"F8", x"E5", x"CD", -- 0x3130,
      x"38", x"44", x"F1", x"F1", x"DD", x"75", x"FC", x"DD", -- 0x3138,
      x"74", x"FD", x"DD", x"73", x"FE", x"DD", x"72", x"FF", -- 0x3140,
      x"D1", x"C1", x"D5", x"C5", x"DD", x"5E", x"FA", x"DD", -- 0x3148,
      x"56", x"FB", x"21", x"35", x"00", x"39", x"01", x"04", -- 0x3150,
      x"00", x"ED", x"B0", x"C1", x"D1", x"21", x"0A", x"00", -- 0x3158,
      x"09", x"DD", x"75", x"FA", x"DD", x"74", x"FB", x"EB", -- 0x3160,
      x"5E", x"23", x"56", x"21", x"1C", x"00", x"19", x"C5", -- 0x3168,
      x"E5", x"CD", x"19", x"36", x"F1", x"DD", x"75", x"FC", -- 0x3170,
      x"DD", x"74", x"FD", x"DD", x"73", x"FE", x"DD", x"72", -- 0x3178,
      x"FF", x"DD", x"5E", x"FA", x"DD", x"56", x"FB", x"21", -- 0x3180,
      x"33", x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", -- 0x3188,
      x"C1", x"69", x"60", x"DD", x"7E", x"F7", x"77", x"23", -- 0x3190,
      x"DD", x"7E", x"F8", x"77", x"21", x"02", x"00", x"09", -- 0x3198,
      x"DD", x"75", x"FE", x"DD", x"74", x"FF", x"DD", x"6E", -- 0x31A0,
      x"F7", x"DD", x"66", x"F8", x"11", x"04", x"00", x"19", -- 0x31A8,
      x"5E", x"23", x"56", x"DD", x"6E", x"FE", x"DD", x"66", -- 0x31B0,
      x"FF", x"73", x"23", x"72", x"21", x"0E", x"00", x"09", -- 0x31B8,
      x"36", x"01", x"21", x"0F", x"00", x"09", x"36", x"00", -- 0x31C0,
      x"21", x"18", x"00", x"09", x"AF", x"77", x"23", x"77", -- 0x31C8,
      x"23", x"77", x"23", x"77", x"21", x"10", x"00", x"09", -- 0x31D0,
      x"AF", x"77", x"23", x"77", x"23", x"77", x"23", x"77", -- 0x31D8,
      x"DD", x"7E", x"F9", x"B7", x"28", x"04", x"AF", x"02", -- 0x31E0,
      x"03", x"02", x"DD", x"6E", x"F9", x"DD", x"F9", x"DD", -- 0x31E8,
      x"E1", x"C9", x"CD", x"13", x"3F", x"2A", x"3F", x"72", -- 0x31F0,
      x"4D", x"7C", x"47", x"B5", x"28", x"02", x"AF", x"02", -- 0x31F8,
      x"DD", x"7E", x"05", x"DD", x"B6", x"04", x"28", x"08", -- 0x3200,
      x"DD", x"4E", x"04", x"DD", x"46", x"05", x"AF", x"02", -- 0x3208,
      x"21", x"3F", x"72", x"DD", x"7E", x"04", x"77", x"23", -- 0x3210,
      x"DD", x"7E", x"05", x"77", x"DD", x"7E", x"08", x"B7", -- 0x3218,
      x"20", x"03", x"6F", x"18", x"09", x"21", x"04", x"00", -- 0x3220,
      x"39", x"E5", x"CD", x"20", x"38", x"F1", x"DD", x"E1", -- 0x3228,
      x"C9", x"CD", x"13", x"3F", x"21", x"F3", x"FF", x"39", -- 0x3230,
      x"F9", x"DD", x"7E", x"04", x"CB", x"7F", x"28", x"1D", -- 0x3238,
      x"E6", x"7F", x"DD", x"77", x"04", x"21", x"00", x"00", -- 0x3240,
      x"E5", x"21", x"00", x"00", x"E5", x"3E", x"37", x"F5", -- 0x3248,
      x"33", x"CD", x"31", x"32", x"F1", x"F1", x"33", x"3E", -- 0x3250,
      x"01", x"95", x"DA", x"49", x"33", x"DD", x"7E", x"04", -- 0x3258,
      x"D6", x"0C", x"3E", x"01", x"28", x"01", x"AF", x"4F", -- 0x3260,
      x"CB", x"41", x"20", x"11", x"C5", x"CD", x"8F", x"35", -- 0x3268,
      x"CD", x"4E", x"33", x"C1", x"7C", x"B5", x"20", x"05", -- 0x3270,
      x"2E", x"FF", x"C3", x"49", x"33", x"21", x"01", x"00", -- 0x3278,
      x"39", x"DD", x"75", x"FA", x"DD", x"74", x"FB", x"DD", -- 0x3280,
      x"46", x"04", x"78", x"CB", x"F7", x"DD", x"6E", x"FA", -- 0x3288,
      x"DD", x"66", x"FB", x"77", x"DD", x"5E", x"FA", x"DD", -- 0x3290,
      x"56", x"FB", x"13", x"DD", x"7E", x"08", x"DD", x"77", -- 0x3298,
      x"FC", x"AF", x"DD", x"77", x"FD", x"DD", x"77", x"FE", -- 0x32A0,
      x"DD", x"77", x"FF", x"DD", x"7E", x"FC", x"12", x"DD", -- 0x32A8,
      x"5E", x"FA", x"DD", x"56", x"FB", x"13", x"13", x"DD", -- 0x32B0,
      x"7E", x"07", x"DD", x"77", x"FC", x"DD", x"7E", x"08", -- 0x32B8,
      x"DD", x"77", x"FD", x"AF", x"DD", x"77", x"FE", x"DD", -- 0x32C0,
      x"77", x"FF", x"DD", x"7E", x"FC", x"12", x"DD", x"6E", -- 0x32C8,
      x"FA", x"DD", x"66", x"FB", x"23", x"23", x"23", x"DD", -- 0x32D0,
      x"5E", x"06", x"73", x"DD", x"7E", x"FA", x"C6", x"04", -- 0x32D8,
      x"5F", x"DD", x"7E", x"FB", x"CE", x"00", x"57", x"DD", -- 0x32E0,
      x"7E", x"05", x"12", x"1E", x"01", x"78", x"B7", x"20", -- 0x32E8,
      x"02", x"1E", x"95", x"DD", x"7E", x"04", x"D6", x"08", -- 0x32F0,
      x"20", x"02", x"1E", x"87", x"DD", x"7E", x"FA", x"C6", -- 0x32F8,
      x"05", x"6F", x"DD", x"7E", x"FB", x"CE", x"00", x"67", -- 0x3300,
      x"73", x"DD", x"5E", x"FA", x"DD", x"56", x"FB", x"C5", -- 0x3308,
      x"21", x"06", x"00", x"E5", x"D5", x"CD", x"A1", x"46", -- 0x3310,
      x"F1", x"F1", x"C1", x"79", x"B7", x"28", x"0E", x"21", -- 0x3318,
      x"00", x"00", x"39", x"01", x"01", x"00", x"C5", x"E5", -- 0x3320,
      x"CD", x"1D", x"3F", x"F1", x"F1", x"0E", x"0A", x"21", -- 0x3328,
      x"00", x"00", x"39", x"C5", x"11", x"01", x"00", x"D5", -- 0x3330,
      x"E5", x"CD", x"1D", x"3F", x"F1", x"F1", x"C1", x"DD", -- 0x3338,
      x"6E", x"F3", x"CB", x"7D", x"28", x"03", x"0D", x"20", -- 0x3340,
      x"E6", x"DD", x"F9", x"DD", x"E1", x"C9", x"3B", x"3A", -- 0x3348,
      x"3D", x"72", x"D3", x"56", x"21", x"00", x"00", x"39", -- 0x3350,
      x"01", x"01", x"00", x"C5", x"E5", x"CD", x"1D", x"3F", -- 0x3358,
      x"F1", x"F1", x"CD", x"69", x"4B", x"7C", x"B5", x"28", -- 0x3360,
      x"05", x"21", x"01", x"00", x"18", x"06", x"CD", x"8F", -- 0x3368,
      x"35", x"21", x"00", x"00", x"33", x"C9", x"CD", x"13", -- 0x3370,
      x"3F", x"F5", x"01", x"E8", x"03", x"21", x"00", x"00", -- 0x3378,
      x"39", x"E5", x"FD", x"E1", x"E5", x"C5", x"11", x"01", -- 0x3380,
      x"00", x"D5", x"FD", x"E5", x"CD", x"1D", x"3F", x"F1", -- 0x3388,
      x"F1", x"C1", x"E1", x"7E", x"3C", x"20", x"15", x"E5", -- 0x3390,
      x"C5", x"3E", x"02", x"F5", x"33", x"CD", x"9F", x"17", -- 0x3398,
      x"33", x"C1", x"E1", x"59", x"50", x"1B", x"4B", x"7A", -- 0x33A0,
      x"47", x"B3", x"20", x"D5", x"7E", x"D6", x"FE", x"28", -- 0x33A8,
      x"05", x"21", x"00", x"00", x"18", x"22", x"E5", x"DD", -- 0x33B0,
      x"4E", x"06", x"DD", x"46", x"07", x"C5", x"DD", x"4E", -- 0x33B8,
      x"04", x"DD", x"46", x"05", x"C5", x"CD", x"1D", x"3F", -- 0x33C0,
      x"F1", x"F1", x"E1", x"01", x"02", x"00", x"C5", x"E5", -- 0x33C8,
      x"CD", x"1D", x"3F", x"F1", x"F1", x"21", x"01", x"00", -- 0x33D0,
      x"F1", x"DD", x"E1", x"C9", x"D1", x"C1", x"C5", x"D5", -- 0x33D8,
      x"79", x"D3", x"BF", x"0E", x"00", x"78", x"D3", x"BF", -- 0x33E0,
      x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", -- 0x33E8,
      x"00", x"00", x"DB", x"BE", x"6F", x"C9", x"CD", x"13", -- 0x33F0,
      x"3F", x"F5", x"F5", x"3B", x"21", x"3C", x"72", x"36", -- 0x33F8,
      x"03", x"21", x"3D", x"72", x"36", x"02", x"3E", x"C8", -- 0x3400,
      x"F5", x"33", x"CD", x"9F", x"17", x"33", x"3A", x"3C", -- 0x3408,
      x"72", x"D3", x"56", x"0E", x"0A", x"21", x"00", x"00", -- 0x3410,
      x"39", x"EB", x"D5", x"FD", x"E1", x"C5", x"D5", x"21", -- 0x3418,
      x"01", x"00", x"E5", x"FD", x"E5", x"CD", x"1D", x"3F", -- 0x3420,
      x"F1", x"F1", x"D1", x"C1", x"79", x"3D", x"4F", x"B7", -- 0x3428,
      x"20", x"E8", x"AF", x"DD", x"77", x"FF", x"D5", x"21", -- 0x3430,
      x"00", x"00", x"E5", x"21", x"00", x"00", x"E5", x"AF", -- 0x3438,
      x"F5", x"33", x"CD", x"31", x"32", x"F1", x"F1", x"33", -- 0x3440,
      x"D1", x"2D", x"C2", x"6C", x"35", x"21", x"3C", x"72", -- 0x3448,
      x"36", x"01", x"21", x"3D", x"72", x"36", x"00", x"D5", -- 0x3450,
      x"21", x"00", x"00", x"E5", x"21", x"AA", x"01", x"E5", -- 0x3458,
      x"3E", x"08", x"F5", x"33", x"CD", x"31", x"32", x"F1", -- 0x3460,
      x"F1", x"33", x"D1", x"2D", x"C2", x"FD", x"34", x"4B", -- 0x3468,
      x"42", x"D5", x"21", x"04", x"00", x"E5", x"C5", x"CD", -- 0x3470,
      x"1D", x"3F", x"F1", x"F1", x"D1", x"6B", x"62", x"23", -- 0x3478,
      x"23", x"7E", x"3D", x"C2", x"6C", x"35", x"6B", x"62", -- 0x3480,
      x"23", x"23", x"23", x"7E", x"D6", x"AA", x"C2", x"6C", -- 0x3488,
      x"35", x"01", x"E8", x"03", x"C5", x"D5", x"21", x"00", -- 0x3490,
      x"40", x"E5", x"21", x"00", x"00", x"E5", x"3E", x"A9", -- 0x3498,
      x"F5", x"33", x"CD", x"31", x"32", x"F1", x"F1", x"33", -- 0x34A0,
      x"7D", x"D1", x"C1", x"B7", x"28", x"11", x"C5", x"D5", -- 0x34A8,
      x"3E", x"14", x"F5", x"33", x"CD", x"9F", x"17", x"33", -- 0x34B0,
      x"D1", x"C1", x"0B", x"78", x"B1", x"20", x"D5", x"78", -- 0x34B8,
      x"B1", x"CA", x"6C", x"35", x"D5", x"21", x"00", x"00", -- 0x34C0,
      x"E5", x"21", x"00", x"00", x"E5", x"3E", x"3A", x"F5", -- 0x34C8,
      x"33", x"CD", x"31", x"32", x"F1", x"F1", x"33", x"7D", -- 0x34D0,
      x"D1", x"B7", x"C2", x"6C", x"35", x"4B", x"42", x"D5", -- 0x34D8,
      x"21", x"04", x"00", x"E5", x"C5", x"CD", x"1D", x"3F", -- 0x34E0,
      x"F1", x"F1", x"D1", x"1A", x"CB", x"77", x"28", x"05", -- 0x34E8,
      x"01", x"0C", x"00", x"18", x"03", x"01", x"04", x"00", -- 0x34F0,
      x"DD", x"71", x"FF", x"18", x"6F", x"21", x"00", x"00", -- 0x34F8,
      x"E5", x"21", x"00", x"00", x"E5", x"3E", x"A9", x"F5", -- 0x3500,
      x"33", x"CD", x"31", x"32", x"F1", x"F1", x"33", x"3E", -- 0x3508,
      x"01", x"95", x"38", x"08", x"DD", x"36", x"FF", x"02", -- 0x3510,
      x"06", x"A9", x"18", x"06", x"DD", x"36", x"FF", x"01", -- 0x3518,
      x"06", x"01", x"11", x"E8", x"03", x"C5", x"D5", x"21", -- 0x3520,
      x"00", x"00", x"E5", x"21", x"00", x"00", x"E5", x"C5", -- 0x3528,
      x"33", x"CD", x"31", x"32", x"F1", x"F1", x"33", x"7D", -- 0x3530,
      x"D1", x"C1", x"B7", x"28", x"11", x"C5", x"D5", x"3E", -- 0x3538,
      x"14", x"F5", x"33", x"CD", x"9F", x"17", x"33", x"D1", -- 0x3540,
      x"C1", x"1B", x"7A", x"B3", x"20", x"D7", x"7A", x"B3", -- 0x3548,
      x"28", x"16", x"21", x"00", x"00", x"E5", x"21", x"00", -- 0x3550,
      x"02", x"E5", x"3E", x"10", x"F5", x"33", x"CD", x"31", -- 0x3558,
      x"32", x"F1", x"F1", x"33", x"7D", x"B7", x"28", x"04", -- 0x3560,
      x"AF", x"DD", x"77", x"FF", x"DD", x"7E", x"FF", x"32", -- 0x3568,
      x"3E", x"72", x"DD", x"7E", x"FF", x"B7", x"28", x"05", -- 0x3570,
      x"01", x"00", x"00", x"18", x"03", x"01", x"01", x"00", -- 0x3578,
      x"21", x"5A", x"73", x"71", x"C5", x"CD", x"8F", x"35", -- 0x3580,
      x"C1", x"69", x"DD", x"F9", x"DD", x"E1", x"C9", x"3B", -- 0x3588,
      x"3A", x"3C", x"72", x"D3", x"56", x"21", x"00", x"00", -- 0x3590,
      x"39", x"01", x"01", x"00", x"C5", x"E5", x"CD", x"1D", -- 0x3598,
      x"3F", x"F1", x"F1", x"33", x"C9", x"CD", x"13", x"3F", -- 0x35A0,
      x"F5", x"3B", x"DD", x"36", x"FD", x"09", x"DD", x"5E", -- 0x35A8,
      x"04", x"DD", x"56", x"05", x"DD", x"7E", x"05", x"DD", -- 0x35B0,
      x"B6", x"04", x"28", x"3B", x"6B", x"62", x"4E", x"23", -- 0x35B8,
      x"46", x"78", x"B1", x"28", x"32", x"0A", x"B7", x"28", -- 0x35C0,
      x"2E", x"6B", x"62", x"23", x"23", x"7E", x"DD", x"77", -- 0x35C8,
      x"FE", x"23", x"7E", x"DD", x"77", x"FF", x"69", x"60", -- 0x35D0,
      x"01", x"04", x"00", x"09", x"4E", x"23", x"46", x"DD", -- 0x35D8,
      x"6E", x"FE", x"DD", x"66", x"FF", x"BF", x"ED", x"42", -- 0x35E0,
      x"20", x"0D", x"D5", x"CD", x"8C", x"2F", x"7D", x"D1", -- 0x35E8,
      x"0F", x"38", x"04", x"AF", x"DD", x"77", x"FD", x"DD", -- 0x35F0,
      x"4E", x"06", x"DD", x"46", x"07", x"DD", x"7E", x"FD", -- 0x35F8,
      x"B7", x"20", x"06", x"EB", x"5E", x"23", x"56", x"18", -- 0x3600,
      x"03", x"11", x"00", x"00", x"7B", x"02", x"03", x"7A", -- 0x3608,
      x"02", x"DD", x"6E", x"FD", x"DD", x"F9", x"DD", x"E1", -- 0x3610,
      x"C9", x"CD", x"13", x"3F", x"F5", x"F5", x"DD", x"6E", -- 0x3618,
      x"04", x"DD", x"66", x"05", x"23", x"23", x"23", x"4E", -- 0x3620,
      x"06", x"00", x"1E", x"00", x"DD", x"71", x"FD", x"DD", -- 0x3628,
      x"70", x"FE", x"DD", x"73", x"FF", x"AF", x"DD", x"77", -- 0x3630,
      x"FC", x"DD", x"6E", x"04", x"DD", x"66", x"05", x"23", -- 0x3638,
      x"23", x"4E", x"06", x"00", x"11", x"00", x"00", x"79", -- 0x3640,
      x"DD", x"B6", x"FC", x"4F", x"78", x"DD", x"B6", x"FD", -- 0x3648,
      x"47", x"7B", x"DD", x"B6", x"FE", x"5F", x"7A", x"DD", -- 0x3650,
      x"B6", x"FF", x"DD", x"71", x"FD", x"DD", x"70", x"FE", -- 0x3658,
      x"DD", x"73", x"FF", x"AF", x"DD", x"77", x"FC", x"DD", -- 0x3660,
      x"6E", x"04", x"DD", x"66", x"05", x"23", x"4E", x"06", -- 0x3668,
      x"00", x"11", x"00", x"00", x"79", x"DD", x"B6", x"FC", -- 0x3670,
      x"4F", x"78", x"DD", x"B6", x"FD", x"47", x"7B", x"DD", -- 0x3678,
      x"B6", x"FE", x"5F", x"7A", x"DD", x"B6", x"FF", x"DD", -- 0x3680,
      x"71", x"FD", x"DD", x"70", x"FE", x"DD", x"73", x"FF", -- 0x3688,
      x"AF", x"DD", x"77", x"FC", x"DD", x"6E", x"04", x"DD", -- 0x3690,
      x"66", x"05", x"4E", x"06", x"00", x"11", x"00", x"00", -- 0x3698,
      x"DD", x"7E", x"FC", x"B1", x"6F", x"DD", x"7E", x"FD", -- 0x36A0,
      x"B0", x"67", x"DD", x"7E", x"FE", x"B3", x"5F", x"DD", -- 0x36A8,
      x"7E", x"FF", x"B2", x"57", x"DD", x"F9", x"DD", x"E1", -- 0x36B0,
      x"C9", x"01", x"03", x"05", x"07", x"09", x"0E", x"10", -- 0x36B8,
      x"12", x"14", x"16", x"18", x"1C", x"1E", x"80", x"9A", -- 0x36C0,
      x"45", x"41", x"8E", x"41", x"8F", x"80", x"45", x"45", -- 0x36C8,
      x"45", x"49", x"49", x"49", x"8E", x"8F", x"90", x"92", -- 0x36D0,
      x"92", x"4F", x"99", x"4F", x"55", x"55", x"59", x"99", -- 0x36D8,
      x"9A", x"9B", x"9C", x"9D", x"9E", x"9F", x"41", x"49", -- 0x36E0,
      x"4F", x"55", x"A5", x"A5", x"A6", x"A7", x"A8", x"A9", -- 0x36E8,
      x"AA", x"AB", x"AC", x"AD", x"AE", x"AF", x"B0", x"B1", -- 0x36F0,
      x"B2", x"B3", x"B4", x"B5", x"B6", x"B7", x"B8", x"B9", -- 0x36F8,
      x"BA", x"BB", x"BC", x"BD", x"BE", x"BF", x"C0", x"C1", -- 0x3700,
      x"C2", x"C3", x"C4", x"C5", x"C6", x"C7", x"C8", x"C9", -- 0x3708,
      x"CA", x"CB", x"CC", x"CD", x"CE", x"CF", x"D0", x"D1", -- 0x3710,
      x"D2", x"D3", x"D4", x"D5", x"D6", x"D7", x"D8", x"D9", -- 0x3718,
      x"DA", x"DB", x"DC", x"DD", x"DE", x"DF", x"E0", x"E1", -- 0x3720,
      x"E2", x"E3", x"E4", x"E5", x"E6", x"E7", x"E8", x"E9", -- 0x3728,
      x"EA", x"EB", x"EC", x"ED", x"EE", x"EF", x"F0", x"F1", -- 0x3730,
      x"F2", x"F3", x"F4", x"F5", x"F6", x"F7", x"F8", x"F9", -- 0x3738,
      x"FA", x"FB", x"FC", x"FD", x"FE", x"FF", x"D1", x"C1", -- 0x3740,
      x"C5", x"D5", x"79", x"D3", x"BF", x"78", x"F6", x"40", -- 0x3748,
      x"D3", x"BF", x"21", x"05", x"00", x"39", x"4E", x"23", -- 0x3750,
      x"46", x"59", x"50", x"0B", x"7A", x"B3", x"C8", x"21", -- 0x3758,
      x"04", x"00", x"39", x"7E", x"D3", x"BE", x"18", x"F1", -- 0x3760,
      x"CD", x"13", x"3F", x"F5", x"F5", x"DD", x"7E", x"06", -- 0x3768,
      x"C6", x"FE", x"DD", x"77", x"06", x"DD", x"7E", x"07", -- 0x3770,
      x"CE", x"FF", x"DD", x"77", x"07", x"DD", x"7E", x"08", -- 0x3778,
      x"CE", x"FF", x"DD", x"77", x"08", x"DD", x"7E", x"09", -- 0x3780,
      x"CE", x"FF", x"DD", x"77", x"09", x"DD", x"4E", x"04", -- 0x3788,
      x"DD", x"46", x"05", x"69", x"60", x"11", x"0C", x"00", -- 0x3790,
      x"19", x"5E", x"23", x"56", x"23", x"23", x"7E", x"2B", -- 0x3798,
      x"6E", x"67", x"7B", x"C6", x"FE", x"5F", x"7A", x"CE", -- 0x37A0,
      x"FF", x"57", x"7D", x"CE", x"FF", x"6F", x"7C", x"CE", -- 0x37A8,
      x"FF", x"67", x"DD", x"7E", x"06", x"93", x"DD", x"7E", -- 0x37B0,
      x"07", x"9A", x"DD", x"7E", x"08", x"9D", x"DD", x"7E", -- 0x37B8,
      x"09", x"9C", x"38", x"07", x"21", x"00", x"00", x"5D", -- 0x37C0,
      x"54", x"18", x"50", x"69", x"60", x"11", x"20", x"00", -- 0x37C8,
      x"19", x"7E", x"DD", x"77", x"FC", x"23", x"7E", x"DD", -- 0x37D0,
      x"77", x"FD", x"23", x"7E", x"DD", x"77", x"FE", x"23", -- 0x37D8,
      x"7E", x"DD", x"77", x"FF", x"69", x"60", x"11", x"08", -- 0x37E0,
      x"00", x"19", x"4E", x"23", x"46", x"11", x"00", x"00", -- 0x37E8,
      x"DD", x"6E", x"08", x"DD", x"66", x"09", x"E5", x"DD", -- 0x37F0,
      x"6E", x"06", x"DD", x"66", x"07", x"E5", x"D5", x"C5", -- 0x37F8,
      x"CD", x"89", x"5D", x"F1", x"F1", x"F1", x"F1", x"7D", -- 0x3800,
      x"DD", x"86", x"FC", x"6F", x"7C", x"DD", x"8E", x"FD", -- 0x3808,
      x"67", x"7B", x"DD", x"8E", x"FE", x"5F", x"7A", x"DD", -- 0x3810,
      x"8E", x"FF", x"57", x"DD", x"F9", x"DD", x"E1", x"C9", -- 0x3818,
      x"CD", x"13", x"3F", x"21", x"CD", x"FF", x"39", x"F9", -- 0x3820,
      x"DD", x"4E", x"04", x"DD", x"46", x"05", x"69", x"60", -- 0x3828,
      x"AF", x"77", x"23", x"77", x"21", x"3F", x"72", x"7E", -- 0x3830,
      x"DD", x"77", x"E5", x"23", x"7E", x"DD", x"77", x"E6", -- 0x3838,
      x"DD", x"B6", x"E5", x"20", x"05", x"2E", x"0C", x"C3", -- 0x3840,
      x"0E", x"3F", x"DD", x"7E", x"E5", x"02", x"03", x"DD", -- 0x3848,
      x"7E", x"E6", x"02", x"DD", x"6E", x"E5", x"DD", x"66", -- 0x3850,
      x"E6", x"7E", x"B7", x"28", x"0C", x"CD", x"8C", x"2F", -- 0x3858,
      x"7D", x"0F", x"38", x"05", x"2E", x"00", x"C3", x"0E", -- 0x3860,
      x"3F", x"DD", x"6E", x"E5", x"DD", x"66", x"E6", x"36", -- 0x3868,
      x"00", x"CD", x"F6", x"33", x"7D", x"0F", x"30", x"05", -- 0x3870,
      x"2E", x"03", x"C3", x"0E", x"3F", x"AF", x"DD", x"77", -- 0x3878,
      x"E7", x"DD", x"77", x"E8", x"DD", x"77", x"E9", x"DD", -- 0x3880,
      x"77", x"EA", x"21", x"00", x"00", x"E5", x"21", x"00", -- 0x3888,
      x"00", x"E5", x"DD", x"6E", x"E5", x"DD", x"66", x"E6", -- 0x3890,
      x"E5", x"CD", x"41", x"52", x"F1", x"F1", x"F1", x"DD", -- 0x3898,
      x"75", x"FE", x"7D", x"D6", x"02", x"C2", x"AF", x"39", -- 0x38A0,
      x"DD", x"7E", x"E5", x"C6", x"28", x"DD", x"77", x"F9", -- 0x38A8,
      x"DD", x"7E", x"E6", x"CE", x"00", x"DD", x"77", x"FA", -- 0x38B0,
      x"21", x"08", x"00", x"39", x"DD", x"75", x"FB", x"DD", -- 0x38B8,
      x"74", x"FC", x"AF", x"DD", x"77", x"FF", x"DD", x"5E", -- 0x38C0,
      x"FF", x"16", x"00", x"6B", x"62", x"29", x"29", x"29", -- 0x38C8,
      x"29", x"01", x"BE", x"01", x"09", x"DD", x"4E", x"F9", -- 0x38D0,
      x"DD", x"46", x"FA", x"09", x"4D", x"44", x"EB", x"29", -- 0x38D8,
      x"29", x"DD", x"7E", x"FB", x"85", x"DD", x"77", x"FD", -- 0x38E0,
      x"DD", x"7E", x"FC", x"8C", x"DD", x"77", x"FE", x"69", -- 0x38E8,
      x"60", x"11", x"04", x"00", x"19", x"7E", x"B7", x"28", -- 0x38F0,
      x"0D", x"21", x"08", x"00", x"09", x"E5", x"CD", x"19", -- 0x38F8,
      x"36", x"F1", x"4D", x"44", x"18", x"06", x"01", x"00", -- 0x3900,
      x"00", x"11", x"00", x"00", x"DD", x"6E", x"FD", x"DD", -- 0x3908,
      x"66", x"FE", x"71", x"23", x"70", x"23", x"73", x"23", -- 0x3910,
      x"72", x"DD", x"34", x"FF", x"DD", x"7E", x"FF", x"D6", -- 0x3918,
      x"04", x"38", x"A3", x"AF", x"DD", x"77", x"FF", x"DD", -- 0x3920,
      x"7E", x"FF", x"DD", x"77", x"FD", x"AF", x"DD", x"77", -- 0x3928,
      x"FE", x"DD", x"7E", x"FD", x"DD", x"77", x"F9", x"DD", -- 0x3930,
      x"7E", x"FE", x"DD", x"77", x"FA", x"3E", x"03", x"18", -- 0x3938,
      x"08", x"DD", x"CB", x"F9", x"26", x"DD", x"CB", x"FA", -- 0x3940,
      x"16", x"3D", x"20", x"F5", x"DD", x"7E", x"FB", x"DD", -- 0x3948,
      x"86", x"F9", x"DD", x"77", x"FD", x"DD", x"7E", x"FC", -- 0x3950,
      x"DD", x"8E", x"FA", x"DD", x"77", x"FE", x"DD", x"5E", -- 0x3958,
      x"FD", x"DD", x"56", x"FE", x"21", x"1A", x"00", x"39", -- 0x3960,
      x"EB", x"01", x"04", x"00", x"ED", x"B0", x"DD", x"7E", -- 0x3968,
      x"EA", x"DD", x"B6", x"E9", x"DD", x"B6", x"E8", x"DD", -- 0x3970,
      x"B6", x"E7", x"28", x"1D", x"DD", x"6E", x"E9", x"DD", -- 0x3978,
      x"66", x"EA", x"E5", x"DD", x"6E", x"E7", x"DD", x"66", -- 0x3980,
      x"E8", x"E5", x"DD", x"6E", x"E5", x"DD", x"66", x"E6", -- 0x3988,
      x"E5", x"CD", x"41", x"52", x"F1", x"F1", x"F1", x"18", -- 0x3990,
      x"03", x"21", x"03", x"00", x"DD", x"75", x"FE", x"7D", -- 0x3998,
      x"D6", x"02", x"38", x"0B", x"DD", x"34", x"FF", x"DD", -- 0x39A0,
      x"7E", x"FF", x"D6", x"04", x"DA", x"27", x"39", x"DD", -- 0x39A8,
      x"7E", x"FE", x"D6", x"04", x"20", x"05", x"2E", x"01", -- 0x39B0,
      x"C3", x"0E", x"3F", x"DD", x"7E", x"FE", x"D6", x"02", -- 0x39B8,
      x"38", x"05", x"2E", x"0D", x"C3", x"0E", x"3F", x"DD", -- 0x39C0,
      x"7E", x"E5", x"C6", x"28", x"DD", x"77", x"EB", x"DD", -- 0x39C8,
      x"7E", x"E6", x"CE", x"00", x"DD", x"77", x"EC", x"DD", -- 0x39D0,
      x"5E", x"EB", x"DD", x"56", x"EC", x"DD", x"6E", x"EB", -- 0x39D8,
      x"DD", x"66", x"EC", x"01", x"0C", x"00", x"09", x"46", -- 0x39E0,
      x"0E", x"00", x"EB", x"11", x"0B", x"00", x"19", x"5E", -- 0x39E8,
      x"16", x"00", x"79", x"B3", x"4F", x"78", x"B2", x"47", -- 0x39F0,
      x"79", x"B7", x"20", x"05", x"78", x"D6", x"02", x"28", -- 0x39F8,
      x"05", x"2E", x"0D", x"C3", x"0E", x"3F", x"DD", x"5E", -- 0x3A00,
      x"EB", x"DD", x"56", x"EC", x"DD", x"6E", x"EB", x"DD", -- 0x3A08,
      x"66", x"EC", x"01", x"17", x"00", x"09", x"46", x"0E", -- 0x3A10,
      x"00", x"EB", x"11", x"16", x"00", x"19", x"5E", x"16", -- 0x3A18,
      x"00", x"79", x"B3", x"4F", x"78", x"B2", x"47", x"17", -- 0x3A20,
      x"9F", x"5F", x"57", x"B3", x"B0", x"B1", x"20", x"13", -- 0x3A28,
      x"DD", x"7E", x"EB", x"C6", x"24", x"4F", x"DD", x"7E", -- 0x3A30,
      x"EC", x"CE", x"00", x"47", x"C5", x"CD", x"19", x"36", -- 0x3A38,
      x"F1", x"4D", x"44", x"DD", x"7E", x"E5", x"C6", x"10", -- 0x3A40,
      x"DD", x"77", x"ED", x"DD", x"7E", x"E6", x"CE", x"00", -- 0x3A48,
      x"DD", x"77", x"EE", x"DD", x"6E", x"ED", x"DD", x"66", -- 0x3A50,
      x"EE", x"71", x"23", x"70", x"23", x"73", x"23", x"72", -- 0x3A58,
      x"DD", x"7E", x"E5", x"C6", x"01", x"DD", x"77", x"FE", -- 0x3A60,
      x"DD", x"7E", x"E6", x"CE", x"00", x"DD", x"77", x"FF", -- 0x3A68,
      x"DD", x"6E", x"EB", x"DD", x"66", x"EC", x"C5", x"01", -- 0x3A70,
      x"10", x"00", x"09", x"C1", x"7E", x"DD", x"6E", x"FE", -- 0x3A78,
      x"DD", x"66", x"FF", x"77", x"DD", x"6E", x"FE", x"DD", -- 0x3A80,
      x"66", x"FF", x"6E", x"3D", x"28", x"0A", x"7D", x"D6", -- 0x3A88,
      x"02", x"28", x"05", x"2E", x"0D", x"C3", x"0E", x"3F", -- 0x3A90,
      x"DD", x"75", x"FC", x"AF", x"DD", x"77", x"FD", x"DD", -- 0x3A98,
      x"77", x"FE", x"DD", x"77", x"FF", x"6F", x"67", x"E5", -- 0x3AA0,
      x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"E5", x"D5", -- 0x3AA8,
      x"C5", x"CD", x"89", x"5D", x"F1", x"F1", x"F1", x"F1", -- 0x3AB0,
      x"DD", x"75", x"EF", x"DD", x"74", x"F0", x"DD", x"73", -- 0x3AB8,
      x"F1", x"DD", x"72", x"F2", x"DD", x"7E", x"E5", x"C6", -- 0x3AC0,
      x"08", x"DD", x"77", x"FA", x"DD", x"7E", x"E6", x"CE", -- 0x3AC8,
      x"00", x"DD", x"77", x"FB", x"DD", x"6E", x"EB", x"DD", -- 0x3AD0,
      x"66", x"EC", x"11", x"0D", x"00", x"19", x"5E", x"16", -- 0x3AD8,
      x"00", x"DD", x"6E", x"FA", x"DD", x"66", x"FB", x"73", -- 0x3AE0,
      x"23", x"72", x"DD", x"6E", x"FA", x"DD", x"66", x"FB", -- 0x3AE8,
      x"4E", x"23", x"46", x"7A", x"B3", x"28", x"0B", x"59", -- 0x3AF0,
      x"50", x"1B", x"79", x"A3", x"4F", x"78", x"A2", x"B1", -- 0x3AF8,
      x"28", x"05", x"2E", x"0D", x"C3", x"0E", x"3F", x"DD", -- 0x3B00,
      x"7E", x"E5", x"C6", x"06", x"DD", x"77", x"F3", x"DD", -- 0x3B08,
      x"7E", x"E6", x"CE", x"00", x"DD", x"77", x"F4", x"DD", -- 0x3B10,
      x"5E", x"EB", x"DD", x"56", x"EC", x"DD", x"6E", x"EB", -- 0x3B18,
      x"DD", x"66", x"EC", x"01", x"12", x"00", x"09", x"46", -- 0x3B20,
      x"0E", x"00", x"EB", x"11", x"11", x"00", x"19", x"5E", -- 0x3B28,
      x"16", x"00", x"79", x"B3", x"4F", x"78", x"B2", x"47", -- 0x3B30,
      x"DD", x"6E", x"F3", x"DD", x"66", x"F4", x"71", x"23", -- 0x3B38,
      x"70", x"79", x"E6", x"0F", x"28", x"05", x"2E", x"0D", -- 0x3B40,
      x"C3", x"0E", x"3F", x"DD", x"5E", x"EB", x"DD", x"56", -- 0x3B48,
      x"EC", x"DD", x"6E", x"EB", x"DD", x"66", x"EC", x"01", -- 0x3B50,
      x"14", x"00", x"09", x"46", x"0E", x"00", x"EB", x"11", -- 0x3B58,
      x"13", x"00", x"19", x"5E", x"16", x"00", x"79", x"B3", -- 0x3B60,
      x"4F", x"78", x"B2", x"47", x"DD", x"71", x"CD", x"78", -- 0x3B68,
      x"DD", x"77", x"CE", x"17", x"9F", x"DD", x"77", x"CF", -- 0x3B70,
      x"DD", x"77", x"D0", x"DD", x"B6", x"CF", x"DD", x"B6", -- 0x3B78,
      x"CE", x"DD", x"B6", x"CD", x"20", x"35", x"DD", x"7E", -- 0x3B80,
      x"EB", x"C6", x"20", x"DD", x"77", x"FE", x"DD", x"7E", -- 0x3B88,
      x"EC", x"CE", x"00", x"DD", x"77", x"FF", x"DD", x"6E", -- 0x3B90,
      x"FE", x"DD", x"66", x"FF", x"E5", x"CD", x"19", x"36", -- 0x3B98,
      x"F1", x"DD", x"75", x"FC", x"DD", x"74", x"FD", x"DD", -- 0x3BA0,
      x"73", x"FE", x"DD", x"72", x"FF", x"21", x"00", x"00", -- 0x3BA8,
      x"39", x"EB", x"21", x"2F", x"00", x"39", x"01", x"04", -- 0x3BB0,
      x"00", x"ED", x"B0", x"DD", x"5E", x"EB", x"DD", x"56", -- 0x3BB8,
      x"EC", x"DD", x"6E", x"EB", x"DD", x"66", x"EC", x"01", -- 0x3BC0,
      x"0F", x"00", x"09", x"46", x"0E", x"00", x"EB", x"11", -- 0x3BC8,
      x"0E", x"00", x"19", x"5E", x"16", x"00", x"79", x"B3", -- 0x3BD0,
      x"5F", x"78", x"B2", x"57", x"4B", x"7A", x"47", x"B3", -- 0x3BD8,
      x"20", x"05", x"2E", x"0D", x"C3", x"0E", x"3F", x"DD", -- 0x3BE0,
      x"71", x"D1", x"DD", x"70", x"D2", x"AF", x"DD", x"77", -- 0x3BE8,
      x"D3", x"DD", x"77", x"D4", x"DD", x"7E", x"D1", x"DD", -- 0x3BF0,
      x"86", x"EF", x"DD", x"77", x"FC", x"DD", x"7E", x"D2", -- 0x3BF8,
      x"DD", x"8E", x"F0", x"DD", x"77", x"FD", x"DD", x"7E", -- 0x3C00,
      x"D3", x"DD", x"8E", x"F1", x"DD", x"77", x"FE", x"DD", -- 0x3C08,
      x"7E", x"D4", x"DD", x"8E", x"F2", x"DD", x"77", x"FF", -- 0x3C10,
      x"DD", x"6E", x"F3", x"DD", x"66", x"F4", x"5E", x"23", -- 0x3C18,
      x"56", x"06", x"04", x"CB", x"3A", x"CB", x"1B", x"10", -- 0x3C20,
      x"FA", x"21", x"00", x"00", x"DD", x"7E", x"FC", x"83", -- 0x3C28,
      x"4F", x"DD", x"7E", x"FD", x"8A", x"47", x"DD", x"7E", -- 0x3C30,
      x"FE", x"8D", x"5F", x"DD", x"7E", x"FF", x"8C", x"57", -- 0x3C38,
      x"DD", x"71", x"F5", x"DD", x"70", x"F6", x"DD", x"73", -- 0x3C40,
      x"F7", x"DD", x"72", x"F8", x"DD", x"7E", x"CD", x"DD", -- 0x3C48,
      x"96", x"F5", x"DD", x"7E", x"CE", x"DD", x"9E", x"F6", -- 0x3C50,
      x"DD", x"7E", x"CF", x"DD", x"9E", x"F7", x"DD", x"7E", -- 0x3C58,
      x"D0", x"DD", x"9E", x"F8", x"30", x"05", x"2E", x"0D", -- 0x3C60,
      x"C3", x"0E", x"3F", x"DD", x"7E", x"CD", x"DD", x"96", -- 0x3C68,
      x"F5", x"DD", x"77", x"FC", x"DD", x"7E", x"CE", x"DD", -- 0x3C70,
      x"9E", x"F6", x"DD", x"77", x"FD", x"DD", x"7E", x"CF", -- 0x3C78,
      x"DD", x"9E", x"F7", x"DD", x"77", x"FE", x"DD", x"7E", -- 0x3C80,
      x"D0", x"DD", x"9E", x"F8", x"DD", x"77", x"FF", x"DD", -- 0x3C88,
      x"6E", x"FA", x"DD", x"66", x"FB", x"4E", x"23", x"46", -- 0x3C90,
      x"11", x"00", x"00", x"D5", x"C5", x"DD", x"6E", x"FE", -- 0x3C98,
      x"DD", x"66", x"FF", x"E5", x"DD", x"6E", x"FC", x"DD", -- 0x3CA0,
      x"66", x"FD", x"E5", x"CD", x"07", x"5F", x"F1", x"F1", -- 0x3CA8,
      x"F1", x"F1", x"7A", x"B3", x"B4", x"B5", x"20", x"05", -- 0x3CB0,
      x"2E", x"0D", x"C3", x"0E", x"3F", x"AF", x"DD", x"77", -- 0x3CB8,
      x"F9", x"3E", x"F5", x"BD", x"3E", x"FF", x"9C", x"3E", -- 0x3CC0,
      x"FF", x"9B", x"3E", x"0F", x"9A", x"38", x"04", x"DD", -- 0x3CC8,
      x"36", x"F9", x"03", x"3E", x"F5", x"BD", x"3E", x"FF", -- 0x3CD0,
      x"9C", x"3E", x"00", x"9B", x"3E", x"00", x"9A", x"38", -- 0x3CD8,
      x"04", x"DD", x"36", x"F9", x"02", x"3E", x"F5", x"BD", -- 0x3CE0,
      x"3E", x"0F", x"9C", x"3E", x"00", x"9B", x"3E", x"00", -- 0x3CE8,
      x"9A", x"38", x"04", x"AF", x"DD", x"77", x"F9", x"DD", -- 0x3CF0,
      x"7E", x"F9", x"B7", x"20", x"05", x"2E", x"0D", x"C3", -- 0x3CF8,
      x"0E", x"3F", x"DD", x"7E", x"E5", x"C6", x"0C", x"DD", -- 0x3D00,
      x"77", x"FA", x"DD", x"7E", x"E6", x"CE", x"00", x"DD", -- 0x3D08,
      x"77", x"FB", x"01", x"02", x"00", x"09", x"4D", x"44", -- 0x3D10,
      x"30", x"01", x"13", x"DD", x"6E", x"FA", x"DD", x"66", -- 0x3D18,
      x"FB", x"71", x"23", x"70", x"23", x"73", x"23", x"72", -- 0x3D20,
      x"DD", x"7E", x"E5", x"C6", x"14", x"5F", x"DD", x"7E", -- 0x3D28,
      x"E6", x"CE", x"00", x"57", x"21", x"1A", x"00", x"39", -- 0x3D30,
      x"01", x"04", x"00", x"ED", x"B0", x"DD", x"7E", x"E5", -- 0x3D38,
      x"C6", x"18", x"DD", x"77", x"FC", x"DD", x"7E", x"E6", -- 0x3D40,
      x"CE", x"00", x"DD", x"77", x"FD", x"DD", x"7E", x"D1", -- 0x3D48,
      x"DD", x"86", x"E7", x"4F", x"DD", x"7E", x"D2", x"DD", -- 0x3D50,
      x"8E", x"E8", x"47", x"DD", x"7E", x"D3", x"DD", x"8E", -- 0x3D58,
      x"E9", x"5F", x"DD", x"7E", x"D4", x"DD", x"8E", x"EA", -- 0x3D60,
      x"57", x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"71", -- 0x3D68,
      x"23", x"70", x"23", x"73", x"23", x"72", x"DD", x"7E", -- 0x3D70,
      x"E5", x"C6", x"20", x"DD", x"77", x"FE", x"DD", x"7E", -- 0x3D78,
      x"E6", x"CE", x"00", x"DD", x"77", x"FF", x"DD", x"7E", -- 0x3D80,
      x"E7", x"DD", x"86", x"F5", x"4F", x"DD", x"7E", x"E8", -- 0x3D88,
      x"DD", x"8E", x"F6", x"47", x"DD", x"7E", x"E9", x"DD", -- 0x3D90,
      x"8E", x"F7", x"5F", x"DD", x"7E", x"EA", x"DD", x"8E", -- 0x3D98,
      x"F8", x"57", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", -- 0x3DA0,
      x"71", x"23", x"70", x"23", x"73", x"23", x"72", x"DD", -- 0x3DA8,
      x"7E", x"E5", x"C6", x"1C", x"DD", x"77", x"FE", x"DD", -- 0x3DB0,
      x"7E", x"E6", x"CE", x"00", x"DD", x"77", x"FF", x"DD", -- 0x3DB8,
      x"7E", x"F9", x"D6", x"03", x"20", x"75", x"DD", x"4E", -- 0x3DC0,
      x"EB", x"DD", x"46", x"EC", x"DD", x"6E", x"EB", x"DD", -- 0x3DC8,
      x"66", x"EC", x"11", x"2B", x"00", x"19", x"56", x"1E", -- 0x3DD0,
      x"00", x"69", x"60", x"01", x"2A", x"00", x"09", x"4E", -- 0x3DD8,
      x"06", x"00", x"7B", x"B1", x"4F", x"7A", x"B0", x"B1", -- 0x3DE0,
      x"28", x"05", x"2E", x"0D", x"C3", x"0E", x"3F", x"DD", -- 0x3DE8,
      x"6E", x"F3", x"DD", x"66", x"F4", x"7E", x"23", x"B6", -- 0x3DF0,
      x"28", x"05", x"2E", x"0D", x"C3", x"0E", x"3F", x"DD", -- 0x3DF8,
      x"7E", x"EB", x"C6", x"2C", x"4F", x"DD", x"7E", x"EC", -- 0x3E00,
      x"CE", x"00", x"47", x"C5", x"CD", x"19", x"36", x"F1", -- 0x3E08,
      x"4D", x"44", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", -- 0x3E10,
      x"71", x"23", x"70", x"23", x"73", x"23", x"72", x"DD", -- 0x3E18,
      x"6E", x"FA", x"DD", x"66", x"FB", x"4E", x"23", x"46", -- 0x3E20,
      x"23", x"5E", x"23", x"56", x"3E", x"02", x"CB", x"21", -- 0x3E28,
      x"CB", x"10", x"CB", x"13", x"CB", x"12", x"3D", x"20", -- 0x3E30,
      x"F5", x"18", x"53", x"DD", x"6E", x"F3", x"DD", x"66", -- 0x3E38,
      x"F4", x"7E", x"23", x"B6", x"20", x"05", x"2E", x"0D", -- 0x3E40,
      x"C3", x"0E", x"3F", x"DD", x"6E", x"FC", x"DD", x"66", -- 0x3E48,
      x"FD", x"4E", x"23", x"46", x"23", x"5E", x"23", x"56", -- 0x3E50,
      x"79", x"DD", x"86", x"EF", x"4F", x"78", x"DD", x"8E", -- 0x3E58,
      x"F0", x"47", x"7B", x"DD", x"8E", x"F1", x"5F", x"7A", -- 0x3E60,
      x"DD", x"8E", x"F2", x"57", x"DD", x"6E", x"FE", x"DD", -- 0x3E68,
      x"66", x"FF", x"71", x"23", x"70", x"23", x"73", x"23", -- 0x3E70,
      x"72", x"DD", x"6E", x"FA", x"DD", x"66", x"FB", x"4E", -- 0x3E78,
      x"23", x"46", x"23", x"5E", x"23", x"56", x"CB", x"21", -- 0x3E80,
      x"CB", x"10", x"CB", x"13", x"CB", x"12", x"D5", x"C5", -- 0x3E88,
      x"DD", x"5E", x"ED", x"DD", x"56", x"EE", x"21", x"33", -- 0x3E90,
      x"00", x"39", x"EB", x"01", x"04", x"00", x"ED", x"B0", -- 0x3E98,
      x"C1", x"D1", x"79", x"C6", x"FF", x"6F", x"78", x"CE", -- 0x3EA0,
      x"01", x"67", x"30", x"01", x"13", x"06", x"09", x"CB", -- 0x3EA8,
      x"3A", x"CB", x"1B", x"CB", x"1C", x"CB", x"1D", x"10", -- 0x3EB0,
      x"F6", x"DD", x"7E", x"FC", x"95", x"DD", x"7E", x"FD", -- 0x3EB8,
      x"9C", x"DD", x"7E", x"FE", x"9B", x"DD", x"7E", x"FF", -- 0x3EC0,
      x"9A", x"30", x"04", x"2E", x"0D", x"18", x"3F", x"DD", -- 0x3EC8,
      x"6E", x"E5", x"DD", x"66", x"E6", x"DD", x"7E", x"F9", -- 0x3ED0,
      x"77", x"DD", x"7E", x"E5", x"C6", x"04", x"4F", x"DD", -- 0x3ED8,
      x"7E", x"E6", x"CE", x"00", x"47", x"2A", x"41", x"72", -- 0x3EE0,
      x"23", x"22", x"41", x"72", x"FD", x"21", x"41", x"72", -- 0x3EE8,
      x"FD", x"7E", x"00", x"02", x"03", x"FD", x"7E", x"01", -- 0x3EF0,
      x"02", x"DD", x"7E", x"E5", x"C6", x"0A", x"4F", x"DD", -- 0x3EF8,
      x"7E", x"E6", x"CE", x"00", x"47", x"3E", x"43", x"02", -- 0x3F00,
      x"03", x"3E", x"72", x"02", x"2E", x"00", x"DD", x"F9", -- 0x3F08,
      x"DD", x"E1", x"C9", x"E1", x"DD", x"E5", x"DD", x"21", -- 0x3F10,
      x"00", x"00", x"DD", x"39", x"E9", x"E5", x"C5", x"D5", -- 0x3F18,
      x"F5", x"21", x"0A", x"00", x"39", x"F9", x"E1", x"D1", -- 0x3F20,
      x"0E", x"57", x"14", x"15", x"28", x"07", x"AF", x"47", -- 0x3F28,
      x"ED", x"B2", x"15", x"18", x"F5", x"1C", x"1D", x"28", -- 0x3F30,
      x"03", x"43", x"ED", x"B2", x"21", x"F2", x"FF", x"39", -- 0x3F38,
      x"F9", x"F1", x"D1", x"C1", x"E1", x"C9", x"CD", x"13", -- 0x3F40,
      x"3F", x"21", x"DD", x"FF", x"39", x"F9", x"21", x"00", -- 0x3F48,
      x"00", x"39", x"DD", x"7E", x"04", x"DD", x"77", x"DF", -- 0x3F50,
      x"DD", x"7E", x"05", x"DD", x"77", x"E0", x"E5", x"DD", -- 0x3F58,
      x"6E", x"DF", x"DD", x"66", x"E0", x"E5", x"CD", x"A5", -- 0x3F60,
      x"35", x"F1", x"F1", x"DD", x"75", x"E1", x"DD", x"7E", -- 0x3F68,
      x"DF", x"C6", x"0F", x"DD", x"77", x"E2", x"DD", x"7E", -- 0x3F70,
      x"E0", x"CE", x"00", x"DD", x"77", x"E3", x"DD", x"7E", -- 0x3F78,
      x"E1", x"B7", x"20", x"0A", x"DD", x"6E", x"E2", x"DD", -- 0x3F80,
      x"66", x"E3", x"7E", x"DD", x"77", x"E1", x"DD", x"7E", -- 0x3F88,
      x"E1", x"B7", x"28", x"06", x"DD", x"6E", x"E1", x"C3", -- 0x3F90,
      x"33", x"44", x"DD", x"7E", x"DF", x"DD", x"77", x"E4", -- 0x3F98,
      x"DD", x"7E", x"E0", x"DD", x"77", x"E5", x"C1", x"E1", -- 0x3FA0,
      x"E5", x"C5", x"11", x"0A", x"00", x"19", x"4E", x"23", -- 0x3FA8,
      x"46", x"23", x"5E", x"23", x"56", x"79", x"DD", x"96", -- 0x3FB0,
      x"06", x"78", x"DD", x"9E", x"07", x"7B", x"DD", x"9E", -- 0x3FB8,
      x"08", x"7A", x"DD", x"9E", x"09", x"30", x"0C", x"DD", -- 0x3FC0,
      x"71", x"06", x"DD", x"70", x"07", x"DD", x"73", x"08", -- 0x3FC8,
      x"DD", x"72", x"09", x"DD", x"7E", x"DF", x"C6", x"10", -- 0x3FD0,
      x"DD", x"77", x"E6", x"DD", x"7E", x"E0", x"CE", x"00", -- 0x3FD8,
      x"DD", x"77", x"E7", x"DD", x"7E", x"E6", x"DD", x"77", -- 0x3FE0,
      x"E8", x"DD", x"7E", x"E7", x"DD", x"77", x"E9", x"DD", -- 0x3FE8,
      x"5E", x"E6", x"DD", x"56", x"E7", x"21", x"0D", x"00", -- 0x3FF0,
      x"39", x"EB", x"01", x"04", x"00", x"ED", x"B0", x"AF", -- 0x3FF8,
      x"DD", x"77", x"EE", x"DD", x"77", x"EF", x"DD", x"77", -- 0x4000,
      x"F0", x"DD", x"77", x"F1", x"DD", x"6E", x"E6", x"DD", -- 0x4008,
      x"66", x"E7", x"AF", x"77", x"23", x"77", x"23", x"77", -- 0x4010,
      x"23", x"77", x"DD", x"7E", x"09", x"DD", x"B6", x"08", -- 0x4018,
      x"DD", x"B6", x"07", x"DD", x"B6", x"06", x"CA", x"8D", -- 0x4020,
      x"43", x"E1", x"E5", x"11", x"08", x"00", x"19", x"4E", -- 0x4028,
      x"23", x"46", x"1E", x"00", x"DD", x"71", x"F3", x"DD", -- 0x4030,
      x"70", x"F4", x"DD", x"73", x"F5", x"AF", x"DD", x"77", -- 0x4038,
      x"F2", x"DD", x"CB", x"F3", x"26", x"DD", x"CB", x"F4", -- 0x4040,
      x"16", x"DD", x"CB", x"F5", x"16", x"DD", x"7E", x"DF", -- 0x4048,
      x"C6", x"14", x"DD", x"77", x"F6", x"DD", x"7E", x"E0", -- 0x4050,
      x"CE", x"00", x"DD", x"77", x"F7", x"DD", x"7E", x"ED", -- 0x4058,
      x"DD", x"B6", x"EC", x"DD", x"B6", x"EB", x"DD", x"B6", -- 0x4060,
      x"EA", x"CA", x"6D", x"41", x"DD", x"7E", x"06", x"C6", -- 0x4068,
      x"FF", x"4F", x"DD", x"7E", x"07", x"CE", x"FF", x"47", -- 0x4070,
      x"DD", x"7E", x"08", x"CE", x"FF", x"5F", x"DD", x"7E", -- 0x4078,
      x"09", x"CE", x"FF", x"57", x"DD", x"6E", x"F4", x"DD", -- 0x4080,
      x"66", x"F5", x"E5", x"DD", x"6E", x"F2", x"DD", x"66", -- 0x4088,
      x"F3", x"E5", x"D5", x"C5", x"CD", x"07", x"5F", x"F1", -- 0x4090,
      x"F1", x"F1", x"F1", x"DD", x"75", x"F8", x"DD", x"74", -- 0x4098,
      x"F9", x"DD", x"73", x"FA", x"DD", x"72", x"FB", x"DD", -- 0x40A0,
      x"7E", x"EA", x"C6", x"FF", x"DD", x"77", x"FC", x"DD", -- 0x40A8,
      x"7E", x"EB", x"CE", x"FF", x"DD", x"77", x"FD", x"DD", -- 0x40B0,
      x"7E", x"EC", x"CE", x"FF", x"DD", x"77", x"FE", x"DD", -- 0x40B8,
      x"7E", x"ED", x"CE", x"FF", x"DD", x"77", x"FF", x"DD", -- 0x40C0,
      x"6E", x"F4", x"DD", x"66", x"F5", x"E5", x"DD", x"6E", -- 0x40C8,
      x"F2", x"DD", x"66", x"F3", x"E5", x"DD", x"6E", x"FE", -- 0x40D0,
      x"DD", x"66", x"FF", x"E5", x"DD", x"6E", x"FC", x"DD", -- 0x40D8,
      x"66", x"FD", x"E5", x"CD", x"07", x"5F", x"F1", x"F1", -- 0x40E0,
      x"F1", x"F1", x"DD", x"7E", x"F8", x"95", x"DD", x"7E", -- 0x40E8,
      x"F9", x"9C", x"DD", x"7E", x"FA", x"9B", x"DD", x"7E", -- 0x40F0,
      x"FB", x"9A", x"38", x"71", x"DD", x"7E", x"F2", x"C6", -- 0x40F8,
      x"FF", x"4F", x"DD", x"7E", x"F3", x"CE", x"FF", x"47", -- 0x4100,
      x"DD", x"7E", x"F4", x"CE", x"FF", x"5F", x"DD", x"7E", -- 0x4108,
      x"F5", x"CE", x"FF", x"2F", x"67", x"79", x"2F", x"F5", -- 0x4110,
      x"78", x"2F", x"4F", x"7B", x"2F", x"6F", x"F1", x"DD", -- 0x4118,
      x"A6", x"FC", x"5F", x"79", x"DD", x"A6", x"FD", x"57", -- 0x4120,
      x"7D", x"DD", x"A6", x"FE", x"4F", x"7C", x"DD", x"A6", -- 0x4128,
      x"FF", x"47", x"DD", x"6E", x"E6", x"DD", x"66", x"E7", -- 0x4130,
      x"73", x"23", x"72", x"23", x"71", x"23", x"70", x"DD", -- 0x4138,
      x"7E", x"06", x"93", x"DD", x"77", x"06", x"DD", x"7E", -- 0x4140,
      x"07", x"9A", x"DD", x"77", x"07", x"DD", x"7E", x"08", -- 0x4148,
      x"99", x"DD", x"77", x"08", x"DD", x"7E", x"09", x"98", -- 0x4150,
      x"DD", x"77", x"09", x"DD", x"5E", x"F6", x"DD", x"56", -- 0x4158,
      x"F7", x"21", x"1F", x"00", x"39", x"EB", x"01", x"04", -- 0x4160,
      x"00", x"ED", x"B0", x"18", x"2A", x"C1", x"E1", x"E5", -- 0x4168,
      x"C5", x"11", x"06", x"00", x"19", x"7E", x"DD", x"77", -- 0x4170,
      x"FC", x"23", x"7E", x"DD", x"77", x"FD", x"23", x"7E", -- 0x4178,
      x"DD", x"77", x"FE", x"23", x"7E", x"DD", x"77", x"FF", -- 0x4180,
      x"DD", x"5E", x"F6", x"DD", x"56", x"F7", x"21", x"1F", -- 0x4188,
      x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", x"DD", -- 0x4190,
      x"7E", x"FF", x"DD", x"B6", x"FE", x"DD", x"B6", x"FD", -- 0x4198,
      x"DD", x"B6", x"FC", x"CA", x"8D", x"43", x"DD", x"7E", -- 0x41A0,
      x"DF", x"DD", x"77", x"FA", x"DD", x"7E", x"E0", x"DD", -- 0x41A8,
      x"77", x"FB", x"DD", x"7E", x"F2", x"DD", x"96", x"06", -- 0x41B0,
      x"DD", x"7E", x"F3", x"DD", x"9E", x"07", x"DD", x"7E", -- 0x41B8,
      x"F4", x"DD", x"9E", x"08", x"DD", x"7E", x"F5", x"DD", -- 0x41C0,
      x"9E", x"09", x"D2", x"BC", x"42", x"DD", x"7E", x"06", -- 0x41C8,
      x"DD", x"96", x"F2", x"DD", x"77", x"06", x"DD", x"7E", -- 0x41D0,
      x"07", x"DD", x"9E", x"F3", x"DD", x"77", x"07", x"DD", -- 0x41D8,
      x"7E", x"08", x"DD", x"9E", x"F4", x"DD", x"77", x"08", -- 0x41E0,
      x"DD", x"7E", x"09", x"DD", x"9E", x"F5", x"DD", x"77", -- 0x41E8,
      x"09", x"DD", x"6E", x"E8", x"DD", x"66", x"E9", x"4E", -- 0x41F0,
      x"23", x"46", x"23", x"5E", x"23", x"56", x"79", x"DD", -- 0x41F8,
      x"86", x"F2", x"4F", x"78", x"DD", x"8E", x"F3", x"47", -- 0x4200,
      x"7B", x"DD", x"8E", x"F4", x"5F", x"7A", x"DD", x"8E", -- 0x4208,
      x"F5", x"57", x"DD", x"6E", x"E8", x"DD", x"66", x"E9", -- 0x4210,
      x"71", x"23", x"70", x"23", x"73", x"23", x"72", x"DD", -- 0x4218,
      x"6E", x"FE", x"DD", x"66", x"FF", x"E5", x"DD", x"6E", -- 0x4220,
      x"FC", x"DD", x"66", x"FD", x"E5", x"DD", x"6E", x"E4", -- 0x4228,
      x"DD", x"66", x"E5", x"E5", x"CD", x"C1", x"44", x"F1", -- 0x4230,
      x"F1", x"F1", x"DD", x"75", x"FC", x"DD", x"74", x"FD", -- 0x4238,
      x"DD", x"73", x"FE", x"DD", x"72", x"FF", x"DD", x"7E", -- 0x4240,
      x"FC", x"DD", x"A6", x"FD", x"DD", x"A6", x"FE", x"DD", -- 0x4248,
      x"A6", x"FF", x"3C", x"20", x"0D", x"DD", x"6E", x"E2", -- 0x4250,
      x"DD", x"66", x"E3", x"36", x"01", x"2E", x"01", x"C3", -- 0x4258,
      x"33", x"44", x"3E", x"01", x"DD", x"BE", x"FC", x"3E", -- 0x4260,
      x"00", x"DD", x"9E", x"FD", x"3E", x"00", x"DD", x"9E", -- 0x4268,
      x"FE", x"3E", x"00", x"DD", x"9E", x"FF", x"30", x"1F", -- 0x4270,
      x"E1", x"E5", x"11", x"0C", x"00", x"19", x"4E", x"23", -- 0x4278,
      x"46", x"23", x"5E", x"23", x"56", x"DD", x"7E", x"FC", -- 0x4280,
      x"91", x"DD", x"7E", x"FD", x"98", x"DD", x"7E", x"FE", -- 0x4288,
      x"9B", x"DD", x"7E", x"FF", x"9A", x"38", x"0D", x"DD", -- 0x4290,
      x"6E", x"E2", x"DD", x"66", x"E3", x"36", x"02", x"2E", -- 0x4298,
      x"02", x"C3", x"33", x"44", x"DD", x"7E", x"FA", x"C6", -- 0x42A0,
      x"14", x"5F", x"DD", x"7E", x"FB", x"CE", x"00", x"57", -- 0x42A8,
      x"21", x"1F", x"00", x"39", x"01", x"04", x"00", x"ED", -- 0x42B0,
      x"B0", x"C3", x"B2", x"41", x"DD", x"6E", x"E6", x"DD", -- 0x42B8,
      x"66", x"E7", x"4E", x"23", x"46", x"23", x"5E", x"23", -- 0x42C0,
      x"56", x"79", x"DD", x"86", x"06", x"4F", x"78", x"DD", -- 0x42C8,
      x"8E", x"07", x"47", x"7B", x"DD", x"8E", x"08", x"5F", -- 0x42D0,
      x"7A", x"DD", x"8E", x"09", x"57", x"DD", x"6E", x"E6", -- 0x42D8,
      x"DD", x"66", x"E7", x"71", x"23", x"70", x"23", x"73", -- 0x42E0,
      x"23", x"72", x"DD", x"7E", x"06", x"B7", x"20", x"07", -- 0x42E8,
      x"DD", x"CB", x"07", x"46", x"CA", x"8D", x"43", x"DD", -- 0x42F0,
      x"6E", x"FE", x"DD", x"66", x"FF", x"E5", x"DD", x"6E", -- 0x42F8,
      x"FC", x"DD", x"66", x"FD", x"E5", x"DD", x"6E", x"DD", -- 0x4300,
      x"DD", x"66", x"DE", x"E5", x"CD", x"68", x"37", x"F1", -- 0x4308,
      x"F1", x"F1", x"DD", x"75", x"FC", x"DD", x"74", x"FD", -- 0x4310,
      x"DD", x"73", x"FE", x"DD", x"72", x"FF", x"21", x"1B", -- 0x4318,
      x"00", x"39", x"EB", x"21", x"1F", x"00", x"39", x"01", -- 0x4320,
      x"04", x"00", x"ED", x"B0", x"DD", x"7E", x"FB", x"DD", -- 0x4328,
      x"B6", x"FA", x"DD", x"B6", x"F9", x"DD", x"B6", x"F8", -- 0x4330,
      x"20", x"0D", x"DD", x"6E", x"E2", x"DD", x"66", x"E3", -- 0x4338,
      x"36", x"02", x"2E", x"02", x"C3", x"33", x"44", x"DD", -- 0x4340,
      x"7E", x"07", x"DD", x"77", x"FC", x"DD", x"7E", x"08", -- 0x4348,
      x"DD", x"77", x"FD", x"DD", x"7E", x"09", x"DD", x"77", -- 0x4350,
      x"FE", x"AF", x"DD", x"77", x"FF", x"DD", x"CB", x"FE", -- 0x4358,
      x"3E", x"DD", x"CB", x"FD", x"1E", x"DD", x"CB", x"FC", -- 0x4360,
      x"1E", x"DD", x"7E", x"FC", x"DD", x"86", x"F8", x"DD", -- 0x4368,
      x"77", x"EE", x"DD", x"7E", x"FD", x"DD", x"8E", x"F9", -- 0x4370,
      x"DD", x"77", x"EF", x"DD", x"7E", x"FE", x"DD", x"8E", -- 0x4378,
      x"FA", x"DD", x"77", x"F0", x"DD", x"7E", x"FF", x"DD", -- 0x4380,
      x"8E", x"FB", x"DD", x"77", x"F1", x"DD", x"5E", x"E6", -- 0x4388,
      x"DD", x"56", x"E7", x"21", x"1F", x"00", x"39", x"EB", -- 0x4390,
      x"01", x"04", x"00", x"ED", x"B0", x"DD", x"7E", x"FC", -- 0x4398,
      x"B7", x"20", x"07", x"DD", x"CB", x"FD", x"46", x"CA", -- 0x43A0,
      x"30", x"44", x"DD", x"7E", x"DF", x"C6", x"18", x"DD", -- 0x43A8,
      x"77", x"FC", x"DD", x"7E", x"E0", x"CE", x"00", x"DD", -- 0x43B0,
      x"77", x"FD", x"DD", x"6E", x"FC", x"DD", x"66", x"FD", -- 0x43B8,
      x"4E", x"23", x"46", x"23", x"5E", x"23", x"56", x"DD", -- 0x43C0,
      x"7E", x"EE", x"91", x"20", x"11", x"DD", x"7E", x"EF", -- 0x43C8,
      x"90", x"20", x"0B", x"DD", x"6E", x"F0", x"DD", x"66", -- 0x43D0,
      x"F1", x"BF", x"ED", x"52", x"28", x"52", x"DD", x"7E", -- 0x43D8,
      x"DF", x"C6", x"1C", x"DD", x"77", x"FE", x"DD", x"7E", -- 0x43E0,
      x"E0", x"CE", x"00", x"DD", x"77", x"FF", x"21", x"01", -- 0x43E8,
      x"00", x"E5", x"DD", x"6E", x"F0", x"DD", x"66", x"F1", -- 0x43F0,
      x"E5", x"DD", x"6E", x"EE", x"DD", x"66", x"EF", x"E5", -- 0x43F8,
      x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"E5", x"CD", -- 0x4400,
      x"61", x"2E", x"F1", x"F1", x"F1", x"F1", x"DD", x"75", -- 0x4408,
      x"FF", x"7D", x"B7", x"28", x"0C", x"DD", x"6E", x"E2", -- 0x4410,
      x"DD", x"66", x"E3", x"36", x"01", x"2E", x"01", x"18", -- 0x4418,
      x"12", x"DD", x"5E", x"FC", x"DD", x"56", x"FD", x"21", -- 0x4420,
      x"11", x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", -- 0x4428,
      x"DD", x"6E", x"E1", x"DD", x"F9", x"DD", x"E1", x"C9", -- 0x4430,
      x"CD", x"13", x"3F", x"F5", x"F5", x"DD", x"7E", x"06", -- 0x4438,
      x"C6", x"1A", x"5F", x"DD", x"7E", x"07", x"CE", x"00", -- 0x4440,
      x"57", x"6B", x"62", x"23", x"46", x"0E", x"00", x"1A", -- 0x4448,
      x"5F", x"16", x"00", x"79", x"B3", x"4F", x"78", x"B2", -- 0x4450,
      x"47", x"DD", x"71", x"FC", x"78", x"DD", x"77", x"FD", -- 0x4458,
      x"17", x"9F", x"DD", x"77", x"FE", x"DD", x"77", x"FF", -- 0x4460,
      x"DD", x"4E", x"04", x"DD", x"46", x"05", x"0A", x"D6", -- 0x4468,
      x"03", x"20", x"3D", x"DD", x"7E", x"06", x"C6", x"14", -- 0x4470,
      x"5F", x"DD", x"7E", x"07", x"CE", x"00", x"57", x"6B", -- 0x4478,
      x"62", x"23", x"46", x"0E", x"00", x"1A", x"5F", x"16", -- 0x4480,
      x"00", x"79", x"B3", x"5F", x"78", x"B2", x"57", x"17", -- 0x4488,
      x"9F", x"01", x"00", x"00", x"DD", x"7E", x"FC", x"B1", -- 0x4490,
      x"DD", x"77", x"FC", x"DD", x"7E", x"FD", x"B0", x"DD", -- 0x4498,
      x"77", x"FD", x"DD", x"7E", x"FE", x"B3", x"DD", x"77", -- 0x44A0,
      x"FE", x"DD", x"7E", x"FF", x"B2", x"DD", x"77", x"FF", -- 0x44A8,
      x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"DD", x"5E", -- 0x44B0,
      x"FE", x"DD", x"56", x"FF", x"DD", x"F9", x"DD", x"E1", -- 0x44B8,
      x"C9", x"CD", x"13", x"3F", x"F5", x"F5", x"F5", x"F5", -- 0x44C0,
      x"DD", x"6E", x"04", x"DD", x"66", x"05", x"4E", x"23", -- 0x44C8,
      x"46", x"DD", x"7E", x"06", x"D6", x"02", x"DD", x"7E", -- 0x44D0,
      x"07", x"DE", x"00", x"DD", x"7E", x"08", x"DE", x"00", -- 0x44D8,
      x"DD", x"7E", x"09", x"DE", x"00", x"38", x"21", x"69", -- 0x44E0,
      x"60", x"11", x"0C", x"00", x"19", x"5E", x"23", x"56", -- 0x44E8,
      x"23", x"23", x"7E", x"2B", x"6E", x"67", x"DD", x"7E", -- 0x44F0,
      x"06", x"93", x"DD", x"7E", x"07", x"9A", x"DD", x"7E", -- 0x44F8,
      x"08", x"9D", x"DD", x"7E", x"09", x"9C", x"38", x"11", -- 0x4500,
      x"DD", x"36", x"F8", x"01", x"AF", x"DD", x"77", x"F9", -- 0x4508,
      x"DD", x"77", x"FA", x"DD", x"77", x"FB", x"C3", x"44", -- 0x4510,
      x"46", x"DD", x"36", x"F8", x"FF", x"DD", x"36", x"F9", -- 0x4518,
      x"FF", x"DD", x"36", x"FA", x"FF", x"DD", x"36", x"FB", -- 0x4520,
      x"FF", x"0A", x"6F", x"79", x"C6", x"18", x"5F", x"78", -- 0x4528,
      x"CE", x"00", x"57", x"7D", x"FE", x"02", x"28", x"07", -- 0x4530,
      x"D6", x"03", x"28", x"7C", x"C3", x"36", x"46", x"C5", -- 0x4538,
      x"21", x"06", x"00", x"39", x"EB", x"01", x"04", x"00", -- 0x4540,
      x"ED", x"B0", x"C1", x"DD", x"5E", x"07", x"DD", x"56", -- 0x4548,
      x"08", x"DD", x"6E", x"09", x"26", x"00", x"DD", x"7E", -- 0x4550,
      x"FC", x"83", x"5F", x"DD", x"7E", x"FD", x"8A", x"57", -- 0x4558,
      x"DD", x"7E", x"FE", x"8D", x"6F", x"DD", x"7E", x"FF", -- 0x4560,
      x"8C", x"67", x"C5", x"E5", x"D5", x"C5", x"CD", x"A2", -- 0x4568,
      x"4D", x"F1", x"F1", x"F1", x"7D", x"C1", x"B7", x"C2", -- 0x4570,
      x"44", x"46", x"21", x"28", x"00", x"09", x"EB", x"DD", -- 0x4578,
      x"6E", x"06", x"DD", x"66", x"07", x"DD", x"4E", x"08", -- 0x4580,
      x"DD", x"46", x"09", x"29", x"CB", x"11", x"CB", x"10", -- 0x4588,
      x"7C", x"E6", x"01", x"67", x"19", x"EB", x"6B", x"62", -- 0x4590,
      x"23", x"46", x"0E", x"00", x"1A", x"5F", x"16", x"00", -- 0x4598,
      x"79", x"B3", x"4F", x"78", x"B2", x"47", x"DD", x"71", -- 0x45A0,
      x"F8", x"78", x"DD", x"77", x"F9", x"17", x"9F", x"DD", -- 0x45A8,
      x"77", x"FA", x"DD", x"77", x"FB", x"C3", x"44", x"46", -- 0x45B0,
      x"C5", x"21", x"06", x"00", x"39", x"EB", x"01", x"04", -- 0x45B8,
      x"00", x"ED", x"B0", x"C1", x"DD", x"5E", x"06", x"DD", -- 0x45C0,
      x"56", x"07", x"DD", x"6E", x"08", x"DD", x"66", x"09", -- 0x45C8,
      x"3E", x"07", x"CB", x"3C", x"CB", x"1D", x"CB", x"1A", -- 0x45D0,
      x"CB", x"1B", x"3D", x"20", x"F5", x"DD", x"7E", x"FC", -- 0x45D8,
      x"83", x"5F", x"DD", x"7E", x"FD", x"8A", x"57", x"DD", -- 0x45E0,
      x"7E", x"FE", x"8D", x"6F", x"DD", x"7E", x"FF", x"8C", -- 0x45E8,
      x"67", x"C5", x"E5", x"D5", x"C5", x"CD", x"A2", x"4D", -- 0x45F0,
      x"F1", x"F1", x"F1", x"7D", x"C1", x"B7", x"20", x"44", -- 0x45F8,
      x"21", x"28", x"00", x"09", x"EB", x"DD", x"6E", x"06", -- 0x4600,
      x"DD", x"66", x"07", x"DD", x"4E", x"08", x"DD", x"46", -- 0x4608,
      x"09", x"3E", x"02", x"29", x"CB", x"11", x"CB", x"10", -- 0x4610,
      x"3D", x"20", x"F8", x"7C", x"E6", x"01", x"67", x"19", -- 0x4618,
      x"E5", x"CD", x"19", x"36", x"F1", x"DD", x"75", x"F8", -- 0x4620,
      x"DD", x"74", x"F9", x"DD", x"73", x"FA", x"7A", x"E6", -- 0x4628,
      x"0F", x"DD", x"77", x"FB", x"18", x"0E", x"DD", x"36", -- 0x4630,
      x"F8", x"01", x"AF", x"DD", x"77", x"F9", x"DD", x"77", -- 0x4638,
      x"FA", x"DD", x"77", x"FB", x"DD", x"6E", x"F8", x"DD", -- 0x4640,
      x"66", x"F9", x"DD", x"5E", x"FA", x"DD", x"56", x"FB", -- 0x4648,
      x"DD", x"F9", x"DD", x"E1", x"C9", x"F5", x"21", x"00", -- 0x4650,
      x"00", x"39", x"FD", x"21", x"04", x"00", x"FD", x"39", -- 0x4658,
      x"FD", x"4E", x"00", x"FD", x"46", x"01", x"C5", x"E5", -- 0x4660,
      x"C5", x"CD", x"A5", x"35", x"F1", x"F1", x"7D", x"C1", -- 0x4668,
      x"5F", x"B7", x"20", x"04", x"AF", x"02", x"03", x"02", -- 0x4670,
      x"6B", x"F1", x"C9", x"F5", x"21", x"00", x"00", x"39", -- 0x4678,
      x"FD", x"21", x"04", x"00", x"FD", x"39", x"FD", x"4E", -- 0x4680,
      x"00", x"FD", x"46", x"01", x"C5", x"E5", x"C5", x"CD", -- 0x4688,
      x"A5", x"35", x"F1", x"F1", x"7D", x"C1", x"5F", x"B7", -- 0x4690,
      x"20", x"04", x"AF", x"02", x"03", x"02", x"6B", x"F1", -- 0x4698,
      x"C9", x"D1", x"C1", x"C5", x"D5", x"21", x"04", x"00", -- 0x46A0,
      x"39", x"5E", x"23", x"56", x"0A", x"D3", x"57", x"03", -- 0x46A8,
      x"1B", x"7A", x"B3", x"20", x"F7", x"C9", x"CD", x"13", -- 0x46B0,
      x"3F", x"21", x"EC", x"FF", x"39", x"F9", x"DD", x"7E", -- 0x46B8,
      x"04", x"DD", x"77", x"F0", x"DD", x"7E", x"05", x"DD", -- 0x46C0,
      x"77", x"F1", x"DD", x"7E", x"F0", x"DD", x"77", x"F2", -- 0x46C8,
      x"DD", x"7E", x"F1", x"DD", x"77", x"F3", x"DD", x"6E", -- 0x46D0,
      x"F0", x"DD", x"66", x"F1", x"7E", x"DD", x"77", x"F4", -- 0x46D8,
      x"23", x"7E", x"DD", x"77", x"F5", x"DD", x"7E", x"08", -- 0x46E0,
      x"D6", x"20", x"DD", x"7E", x"09", x"DE", x"00", x"30", -- 0x46E8,
      x"07", x"DD", x"7E", x"06", x"E6", x"1F", x"28", x"05", -- 0x46F0,
      x"2E", x"02", x"C3", x"C5", x"49", x"DD", x"7E", x"F0", -- 0x46F8,
      x"C6", x"0E", x"5F", x"DD", x"7E", x"F1", x"CE", x"00", -- 0x4700,
      x"57", x"21", x"1A", x"00", x"39", x"01", x"04", x"00", -- 0x4708,
      x"ED", x"B0", x"DD", x"6E", x"F0", x"DD", x"66", x"F1", -- 0x4710,
      x"11", x"06", x"00", x"19", x"7E", x"DD", x"77", x"F6", -- 0x4718,
      x"23", x"7E", x"DD", x"77", x"F7", x"23", x"7E", x"DD", -- 0x4720,
      x"77", x"F8", x"23", x"7E", x"DD", x"77", x"F9", x"DD", -- 0x4728,
      x"7E", x"F4", x"C6", x"1C", x"DD", x"77", x"FE", x"DD", -- 0x4730,
      x"7E", x"F5", x"CE", x"00", x"DD", x"77", x"FF", x"DD", -- 0x4738,
      x"7E", x"F9", x"DD", x"B6", x"F8", x"DD", x"B6", x"F7", -- 0x4740,
      x"DD", x"B6", x"F6", x"20", x"1B", x"DD", x"6E", x"F4", -- 0x4748,
      x"DD", x"66", x"F5", x"7E", x"D6", x"03", x"38", x"10", -- 0x4750,
      x"DD", x"5E", x"FE", x"DD", x"56", x"FF", x"21", x"0A", -- 0x4758,
      x"00", x"39", x"EB", x"01", x"04", x"00", x"ED", x"B0", -- 0x4760,
      x"DD", x"7E", x"F0", x"C6", x"16", x"DD", x"77", x"FA", -- 0x4768,
      x"DD", x"7E", x"F1", x"CE", x"00", x"DD", x"77", x"FB", -- 0x4770,
      x"DD", x"7E", x"F9", x"DD", x"B6", x"F8", x"DD", x"B6", -- 0x4778,
      x"F7", x"DD", x"B6", x"F6", x"20", x"69", x"DD", x"4E", -- 0x4780,
      x"06", x"DD", x"46", x"07", x"DD", x"5E", x"08", x"DD", -- 0x4788,
      x"56", x"09", x"3E", x"05", x"CB", x"3A", x"CB", x"1B", -- 0x4790,
      x"CB", x"18", x"CB", x"19", x"3D", x"20", x"F5", x"DD", -- 0x4798,
      x"6E", x"F4", x"DD", x"66", x"F5", x"C5", x"01", x"06", -- 0x47A0,
      x"00", x"09", x"C1", x"7E", x"23", x"66", x"DD", x"77", -- 0x47A8,
      x"EC", x"DD", x"74", x"ED", x"AF", x"DD", x"77", x"EE", -- 0x47B0,
      x"DD", x"77", x"EF", x"79", x"DD", x"96", x"EC", x"78", -- 0x47B8,
      x"DD", x"9E", x"ED", x"7B", x"DD", x"9E", x"EE", x"7A", -- 0x47C0,
      x"DD", x"9E", x"EF", x"38", x"05", x"2E", x"02", x"C3", -- 0x47C8,
      x"C5", x"49", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", -- 0x47D0,
      x"4E", x"23", x"46", x"23", x"5E", x"23", x"56", x"DD", -- 0x47D8,
      x"6E", x"FA", x"DD", x"66", x"FB", x"71", x"23", x"70", -- 0x47E0,
      x"23", x"73", x"23", x"72", x"C3", x"02", x"49", x"DD", -- 0x47E8,
      x"6E", x"F4", x"DD", x"66", x"F5", x"11", x"08", x"00", -- 0x47F0,
      x"19", x"4E", x"23", x"46", x"1E", x"00", x"DD", x"71", -- 0x47F8,
      x"FD", x"DD", x"70", x"FE", x"DD", x"73", x"FF", x"AF", -- 0x4800,
      x"DD", x"77", x"FC", x"DD", x"CB", x"FD", x"26", x"DD", -- 0x4808,
      x"CB", x"FE", x"16", x"DD", x"CB", x"FF", x"16", x"DD", -- 0x4810,
      x"4E", x"F4", x"DD", x"46", x"F5", x"DD", x"7E", x"06", -- 0x4818,
      x"DD", x"96", x"FC", x"DD", x"7E", x"07", x"DD", x"9E", -- 0x4820,
      x"FD", x"DD", x"7E", x"08", x"DD", x"9E", x"FE", x"DD", -- 0x4828,
      x"7E", x"09", x"DD", x"9E", x"FF", x"DA", x"D8", x"48", -- 0x4830,
      x"C5", x"DD", x"6E", x"F8", x"DD", x"66", x"F9", x"E5", -- 0x4838,
      x"DD", x"6E", x"F6", x"DD", x"66", x"F7", x"E5", x"DD", -- 0x4840,
      x"6E", x"F2", x"DD", x"66", x"F3", x"E5", x"CD", x"C1", -- 0x4848,
      x"44", x"F1", x"F1", x"F1", x"C1", x"DD", x"75", x"F6", -- 0x4850,
      x"DD", x"74", x"F7", x"DD", x"73", x"F8", x"DD", x"72", -- 0x4858,
      x"F9", x"DD", x"7E", x"F6", x"DD", x"A6", x"F7", x"DD", -- 0x4860,
      x"A6", x"F8", x"DD", x"A6", x"F9", x"3C", x"20", x"05", -- 0x4868,
      x"2E", x"01", x"C3", x"C5", x"49", x"DD", x"7E", x"F6", -- 0x4870,
      x"D6", x"02", x"DD", x"7E", x"F7", x"DE", x"00", x"DD", -- 0x4878,
      x"7E", x"F8", x"DE", x"00", x"DD", x"7E", x"F9", x"DE", -- 0x4880,
      x"00", x"38", x"21", x"69", x"60", x"11", x"0C", x"00", -- 0x4888,
      x"19", x"5E", x"23", x"56", x"23", x"23", x"7E", x"2B", -- 0x4890,
      x"6E", x"67", x"DD", x"7E", x"F6", x"93", x"DD", x"7E", -- 0x4898,
      x"F7", x"9A", x"DD", x"7E", x"F8", x"9D", x"DD", x"7E", -- 0x48A0,
      x"F9", x"9C", x"38", x"05", x"2E", x"02", x"C3", x"C5", -- 0x48A8,
      x"49", x"DD", x"7E", x"06", x"DD", x"96", x"FC", x"DD", -- 0x48B0,
      x"77", x"06", x"DD", x"7E", x"07", x"DD", x"9E", x"FD", -- 0x48B8,
      x"DD", x"77", x"07", x"DD", x"7E", x"08", x"DD", x"9E", -- 0x48C0,
      x"FE", x"DD", x"77", x"08", x"DD", x"7E", x"09", x"DD", -- 0x48C8,
      x"9E", x"FF", x"DD", x"77", x"09", x"C3", x"1D", x"48", -- 0x48D0,
      x"DD", x"6E", x"F8", x"DD", x"66", x"F9", x"E5", x"DD", -- 0x48D8,
      x"6E", x"F6", x"DD", x"66", x"F7", x"E5", x"DD", x"6E", -- 0x48E0,
      x"F4", x"DD", x"66", x"F5", x"E5", x"CD", x"68", x"37", -- 0x48E8,
      x"F1", x"F1", x"F1", x"4D", x"44", x"DD", x"6E", x"FA", -- 0x48F0,
      x"DD", x"66", x"FB", x"71", x"23", x"70", x"23", x"73", -- 0x48F8,
      x"23", x"72", x"DD", x"7E", x"F0", x"C6", x"12", x"5F", -- 0x4900,
      x"DD", x"7E", x"F1", x"CE", x"00", x"57", x"21", x"0A", -- 0x4908,
      x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", x"DD", -- 0x4910,
      x"5E", x"FA", x"DD", x"56", x"FB", x"21", x"10", x"00", -- 0x4918,
      x"39", x"EB", x"01", x"04", x"00", x"ED", x"B0", x"DD", -- 0x4920,
      x"7E", x"FF", x"DD", x"B6", x"FE", x"DD", x"B6", x"FD", -- 0x4928,
      x"DD", x"B6", x"FC", x"20", x"05", x"2E", x"02", x"C3", -- 0x4930,
      x"C5", x"49", x"DD", x"4E", x"07", x"DD", x"46", x"08", -- 0x4938,
      x"DD", x"5E", x"09", x"16", x"00", x"CB", x"3B", x"CB", -- 0x4940,
      x"18", x"CB", x"19", x"79", x"DD", x"86", x"FC", x"4F", -- 0x4948,
      x"78", x"DD", x"8E", x"FD", x"47", x"7B", x"DD", x"8E", -- 0x4950,
      x"FE", x"5F", x"7A", x"DD", x"8E", x"FF", x"57", x"DD", -- 0x4958,
      x"6E", x"FA", x"DD", x"66", x"FB", x"71", x"23", x"70", -- 0x4960,
      x"23", x"73", x"23", x"72", x"DD", x"7E", x"F0", x"C6", -- 0x4968,
      x"1A", x"DD", x"77", x"FE", x"DD", x"7E", x"F1", x"CE", -- 0x4970,
      x"00", x"DD", x"77", x"FF", x"DD", x"7E", x"F4", x"C6", -- 0x4978,
      x"28", x"DD", x"77", x"FC", x"DD", x"7E", x"F5", x"CE", -- 0x4980,
      x"00", x"DD", x"77", x"FD", x"DD", x"7E", x"06", x"DD", -- 0x4988,
      x"77", x"F6", x"DD", x"7E", x"07", x"E6", x"01", x"DD", -- 0x4990,
      x"77", x"F7", x"DD", x"36", x"F8", x"00", x"DD", x"36", -- 0x4998,
      x"F9", x"00", x"DD", x"7E", x"F6", x"DD", x"86", x"FC", -- 0x49A0,
      x"DD", x"77", x"FA", x"DD", x"7E", x"F7", x"DD", x"8E", -- 0x49A8,
      x"FD", x"DD", x"77", x"FB", x"DD", x"6E", x"FE", x"DD", -- 0x49B0,
      x"66", x"FF", x"DD", x"7E", x"FA", x"77", x"23", x"DD", -- 0x49B8,
      x"7E", x"FB", x"77", x"2E", x"00", x"DD", x"F9", x"DD", -- 0x49C0,
      x"E1", x"C9", x"CD", x"13", x"3F", x"21", x"F6", x"FF", -- 0x49C8,
      x"39", x"F9", x"DD", x"7E", x"04", x"DD", x"77", x"F6", -- 0x49D0,
      x"DD", x"7E", x"05", x"DD", x"77", x"F7", x"C1", x"C5", -- 0x49D8,
      x"E1", x"E5", x"7E", x"DD", x"77", x"F8", x"23", x"7E", -- 0x49E0,
      x"DD", x"77", x"F9", x"DD", x"5E", x"06", x"DD", x"56", -- 0x49E8,
      x"07", x"1A", x"D6", x"2F", x"20", x"09", x"13", x"DD", -- 0x49F0,
      x"73", x"06", x"DD", x"72", x"07", x"18", x"F2", x"DD", -- 0x49F8,
      x"73", x"06", x"DD", x"72", x"07", x"21", x"06", x"00", -- 0x4A00,
      x"09", x"AF", x"77", x"23", x"77", x"23", x"77", x"23", -- 0x4A08,
      x"77", x"DD", x"5E", x"06", x"DD", x"56", x"07", x"1A", -- 0x4A10,
      x"5F", x"17", x"9F", x"57", x"7B", x"D6", x"20", x"7A", -- 0x4A18,
      x"DE", x"00", x"30", x"19", x"21", x"27", x"00", x"09", -- 0x4A20,
      x"36", x"80", x"21", x"00", x"00", x"E5", x"21", x"00", -- 0x4A28,
      x"00", x"E5", x"C5", x"CD", x"B6", x"46", x"F1", x"F1", -- 0x4A30,
      x"F1", x"5D", x"C3", x"EE", x"4A", x"21", x"10", x"00", -- 0x4A38,
      x"39", x"C5", x"E5", x"C5", x"CD", x"31", x"4E", x"F1", -- 0x4A40,
      x"F1", x"7D", x"C1", x"5F", x"B7", x"C2", x"EE", x"4A", -- 0x4A48,
      x"C5", x"C5", x"CD", x"54", x"55", x"F1", x"7D", x"C1", -- 0x4A50,
      x"5F", x"E1", x"E5", x"C5", x"01", x"27", x"00", x"09", -- 0x4A58,
      x"C1", x"7E", x"E6", x"04", x"57", x"2E", x"00", x"7B", -- 0x4A60,
      x"B7", x"28", x"0E", x"7B", x"D6", x"04", x"C2", x"EE", -- 0x4A68,
      x"4A", x"7D", x"B2", x"20", x"79", x"1E", x"05", x"18", -- 0x4A70,
      x"75", x"7D", x"B2", x"20", x"71", x"E1", x"E5", x"11", -- 0x4A78,
      x"04", x"00", x"19", x"CB", x"66", x"20", x"04", x"1E", -- 0x4A80,
      x"05", x"18", x"63", x"DD", x"7E", x"F6", x"C6", x"06", -- 0x4A88,
      x"DD", x"77", x"FA", x"DD", x"7E", x"F7", x"CE", x"00", -- 0x4A90,
      x"DD", x"77", x"FB", x"DD", x"7E", x"F8", x"C6", x"28", -- 0x4A98,
      x"DD", x"77", x"FE", x"DD", x"7E", x"F9", x"CE", x"00", -- 0x4AA0,
      x"DD", x"77", x"FF", x"E1", x"E5", x"11", x"0E", x"00", -- 0x4AA8,
      x"19", x"5E", x"23", x"7E", x"E6", x"01", x"57", x"7B", -- 0x4AB0,
      x"DD", x"86", x"FE", x"5F", x"7A", x"DD", x"8E", x"FF", -- 0x4AB8,
      x"57", x"C5", x"D5", x"DD", x"6E", x"F8", x"DD", x"66", -- 0x4AC0,
      x"F9", x"E5", x"CD", x"38", x"44", x"F1", x"F1", x"DD", -- 0x4AC8,
      x"75", x"FC", x"DD", x"74", x"FD", x"DD", x"73", x"FE", -- 0x4AD0,
      x"DD", x"72", x"FF", x"DD", x"5E", x"FA", x"DD", x"56", -- 0x4AD8,
      x"FB", x"21", x"08", x"00", x"39", x"01", x"04", x"00", -- 0x4AE0,
      x"ED", x"B0", x"C1", x"C3", x"3D", x"4A", x"6B", x"DD", -- 0x4AE8,
      x"F9", x"DD", x"E1", x"C9", x"F5", x"21", x"00", x"00", -- 0x4AF0,
      x"39", x"FD", x"21", x"04", x"00", x"FD", x"39", x"FD", -- 0x4AF8,
      x"4E", x"00", x"FD", x"46", x"01", x"C5", x"E5", x"C5", -- 0x4B00,
      x"CD", x"A5", x"35", x"F1", x"F1", x"C1", x"7D", x"B7", -- 0x4B08,
      x"20", x"55", x"21", x"07", x"00", x"39", x"7E", x"2B", -- 0x4B10,
      x"B6", x"20", x"11", x"21", x"00", x"00", x"E5", x"21", -- 0x4B18,
      x"00", x"00", x"E5", x"C5", x"CD", x"B6", x"46", x"F1", -- 0x4B20,
      x"F1", x"F1", x"18", x"3B", x"C5", x"21", x"00", x"00", -- 0x4B28,
      x"E5", x"C5", x"CD", x"2A", x"53", x"F1", x"F1", x"C1", -- 0x4B30,
      x"7D", x"D6", x"04", x"20", x"01", x"6F", x"7D", x"B7", -- 0x4B38,
      x"20", x"25", x"21", x"06", x"00", x"39", x"7E", x"23", -- 0x4B40,
      x"66", x"6F", x"E5", x"C5", x"CD", x"A5", x"4B", x"F1", -- 0x4B48,
      x"21", x"00", x"00", x"E3", x"21", x"06", x"00", x"39", -- 0x4B50,
      x"4E", x"23", x"46", x"C5", x"CD", x"0B", x"59", x"F1", -- 0x4B58,
      x"F1", x"7D", x"D6", x"04", x"20", x"01", x"6F", x"F1", -- 0x4B60,
      x"C9", x"CD", x"13", x"3F", x"3B", x"01", x"88", x"13", -- 0x4B68,
      x"21", x"00", x"00", x"39", x"C5", x"11", x"01", x"00", -- 0x4B70,
      x"D5", x"E5", x"CD", x"1D", x"3F", x"F1", x"F1", x"C1", -- 0x4B78,
      x"DD", x"7E", x"FF", x"3C", x"28", x"0F", x"C5", x"3E", -- 0x4B80,
      x"02", x"F5", x"33", x"CD", x"9F", x"17", x"33", x"C1", -- 0x4B88,
      x"0B", x"78", x"B1", x"20", x"DB", x"78", x"B1", x"28", -- 0x4B90,
      x"05", x"21", x"01", x"00", x"18", x"03", x"21", x"00", -- 0x4B98,
      x"00", x"33", x"DD", x"E1", x"C9", x"CD", x"13", x"3F", -- 0x4BA0,
      x"21", x"EF", x"FF", x"39", x"F9", x"DD", x"7E", x"04", -- 0x4BA8,
      x"DD", x"77", x"EF", x"DD", x"7E", x"05", x"DD", x"77", -- 0x4BB0,
      x"F0", x"E1", x"E5", x"7E", x"DD", x"77", x"FE", x"23", -- 0x4BB8,
      x"7E", x"DD", x"77", x"FF", x"DD", x"7E", x"06", x"DD", -- 0x4BC0,
      x"77", x"F1", x"DD", x"7E", x"07", x"DD", x"77", x"F2", -- 0x4BC8,
      x"DD", x"7E", x"F1", x"C6", x"05", x"DD", x"77", x"F3", -- 0x4BD0,
      x"DD", x"7E", x"F2", x"CE", x"00", x"DD", x"77", x"F4", -- 0x4BD8,
      x"DD", x"6E", x"F3", x"DD", x"66", x"F4", x"36", x"00", -- 0x4BE0,
      x"E1", x"E5", x"11", x"16", x"00", x"19", x"4E", x"23", -- 0x4BE8,
      x"46", x"23", x"7E", x"23", x"B6", x"B0", x"B1", x"CA", -- 0x4BF0,
      x"9D", x"4D", x"E1", x"E5", x"11", x"28", x"00", x"19", -- 0x4BF8,
      x"4E", x"23", x"46", x"23", x"5E", x"23", x"56", x"DD", -- 0x4C00,
      x"7E", x"F1", x"C6", x"05", x"DD", x"77", x"F5", x"DD", -- 0x4C08,
      x"7E", x"F2", x"CE", x"00", x"DD", x"77", x"F6", x"79", -- 0x4C10,
      x"A0", x"A3", x"A2", x"3C", x"CA", x"AB", x"4C", x"AF", -- 0x4C18,
      x"DD", x"77", x"F7", x"0E", x"00", x"DD", x"7E", x"F5", -- 0x4C20,
      x"DD", x"77", x"F8", x"DD", x"7E", x"F6", x"DD", x"77", -- 0x4C28,
      x"F9", x"DD", x"7E", x"FE", x"DD", x"77", x"FA", x"DD", -- 0x4C30,
      x"7E", x"FF", x"DD", x"77", x"FB", x"AF", x"DD", x"77", -- 0x4C38,
      x"FE", x"AF", x"DD", x"77", x"FF", x"DD", x"6E", x"FA", -- 0x4C40,
      x"DD", x"66", x"FB", x"11", x"0A", x"00", x"19", x"5E", -- 0x4C48,
      x"23", x"56", x"DD", x"6E", x"FE", x"26", x"00", x"29", -- 0x4C50,
      x"19", x"7E", x"DD", x"77", x"FC", x"23", x"7E", x"DD", -- 0x4C58,
      x"77", x"FD", x"DD", x"B6", x"FC", x"28", x"31", x"DD", -- 0x4C60,
      x"7E", x"FF", x"D6", x"FE", x"38", x"04", x"0E", x"00", -- 0x4C68,
      x"18", x"26", x"DD", x"34", x"FE", x"DD", x"46", x"FC", -- 0x4C70,
      x"DD", x"5E", x"FF", x"DD", x"34", x"FF", x"DD", x"4E", -- 0x4C78,
      x"FF", x"DD", x"6E", x"F8", x"DD", x"66", x"F9", x"16", -- 0x4C80,
      x"00", x"19", x"78", x"77", x"B7", x"20", x"03", x"4F", -- 0x4C88,
      x"18", x"06", x"AF", x"DD", x"77", x"F7", x"18", x"AD", -- 0x4C90,
      x"DD", x"7E", x"F7", x"B7", x"28", x"02", x"0E", x"00", -- 0x4C98,
      x"DD", x"6E", x"F8", x"DD", x"66", x"F9", x"06", x"00", -- 0x4CA0,
      x"09", x"36", x"00", x"0E", x"00", x"DD", x"6E", x"F3", -- 0x4CA8,
      x"DD", x"66", x"F4", x"46", x"DD", x"7E", x"EF", x"C6", -- 0x4CB0,
      x"1A", x"5F", x"DD", x"7E", x"F0", x"CE", x"00", x"57", -- 0x4CB8,
      x"78", x"B7", x"C2", x"41", x"4D", x"DD", x"73", x"F9", -- 0x4CC0,
      x"DD", x"72", x"FA", x"DD", x"7E", x"F5", x"DD", x"77", -- 0x4CC8,
      x"FB", x"DD", x"7E", x"F6", x"DD", x"77", x"FC", x"DD", -- 0x4CD0,
      x"7E", x"F5", x"DD", x"77", x"FD", x"DD", x"7E", x"F6", -- 0x4CD8,
      x"DD", x"77", x"FE", x"AF", x"DD", x"77", x"FF", x"DD", -- 0x4CE0,
      x"7E", x"FF", x"D6", x"0B", x"30", x"48", x"DD", x"6E", -- 0x4CE8,
      x"F9", x"DD", x"66", x"FA", x"46", x"23", x"66", x"78", -- 0x4CF0,
      x"DD", x"86", x"FF", x"6F", x"30", x"01", x"24", x"DD", -- 0x4CF8,
      x"34", x"FF", x"46", x"78", x"FE", x"20", x"28", x"DF", -- 0x4D00,
      x"D6", x"05", x"20", x"02", x"06", x"E5", x"DD", x"7E", -- 0x4D08,
      x"FF", x"D6", x"09", x"20", x"12", x"79", x"FE", x"0C", -- 0x4D10,
      x"30", x"0D", x"0C", x"DD", x"86", x"FB", x"6F", x"3E", -- 0x4D18,
      x"00", x"DD", x"8E", x"FC", x"67", x"36", x"2E", x"79", -- 0x4D20,
      x"0C", x"DD", x"86", x"FD", x"6F", x"3E", x"00", x"DD", -- 0x4D28,
      x"8E", x"FE", x"67", x"70", x"18", x"B1", x"DD", x"6E", -- 0x4D30,
      x"FB", x"DD", x"66", x"FC", x"06", x"00", x"09", x"36", -- 0x4D38,
      x"00", x"DD", x"6E", x"F3", x"DD", x"66", x"F4", x"7E", -- 0x4D40,
      x"B7", x"20", x"1C", x"B1", x"20", x"0E", x"79", x"0C", -- 0x4D48,
      x"DD", x"86", x"F5", x"6F", x"3E", x"00", x"DD", x"8E", -- 0x4D50,
      x"F6", x"67", x"36", x"3F", x"DD", x"6E", x"F5", x"DD", -- 0x4D58,
      x"66", x"F6", x"06", x"00", x"09", x"36", x"00", x"DD", -- 0x4D60,
      x"7E", x"F1", x"C6", x"04", x"4F", x"DD", x"7E", x"F2", -- 0x4D68,
      x"CE", x"00", x"47", x"6B", x"62", x"7E", x"23", x"66", -- 0x4D70,
      x"6F", x"C5", x"01", x"0B", x"00", x"09", x"C1", x"7E", -- 0x4D78,
      x"02", x"EB", x"4E", x"23", x"46", x"21", x"1C", x"00", -- 0x4D80,
      x"09", x"E5", x"CD", x"19", x"36", x"F1", x"4D", x"44", -- 0x4D88,
      x"DD", x"6E", x"F1", x"DD", x"66", x"F2", x"71", x"23", -- 0x4D90,
      x"70", x"23", x"73", x"23", x"72", x"DD", x"F9", x"DD", -- 0x4D98,
      x"E1", x"C9", x"CD", x"13", x"3F", x"F5", x"F5", x"3B", -- 0x4DA0,
      x"AF", x"DD", x"77", x"FB", x"DD", x"4E", x"04", x"DD", -- 0x4DA8,
      x"46", x"05", x"21", x"24", x"00", x"09", x"EB", x"D5", -- 0x4DB0,
      x"C5", x"21", x"05", x"00", x"39", x"EB", x"01", x"04", -- 0x4DB8,
      x"00", x"ED", x"B0", x"C1", x"D1", x"DD", x"7E", x"06", -- 0x4DC0,
      x"DD", x"96", x"FC", x"20", x"18", x"DD", x"7E", x"07", -- 0x4DC8,
      x"DD", x"96", x"FD", x"20", x"10", x"DD", x"7E", x"08", -- 0x4DD0,
      x"DD", x"96", x"FE", x"20", x"08", x"DD", x"7E", x"09", -- 0x4DD8,
      x"DD", x"96", x"FF", x"28", x"44", x"FD", x"21", x"28", -- 0x4DE0,
      x"00", x"FD", x"09", x"D5", x"21", x"01", x"00", x"E5", -- 0x4DE8,
      x"DD", x"6E", x"08", x"DD", x"66", x"09", x"E5", x"DD", -- 0x4DF0,
      x"6E", x"06", x"DD", x"66", x"07", x"E5", x"FD", x"E5", -- 0x4DF8,
      x"CD", x"61", x"2E", x"F1", x"F1", x"F1", x"F1", x"7D", -- 0x4E00,
      x"D1", x"B7", x"28", x"14", x"DD", x"36", x"06", x"FF", -- 0x4E08,
      x"DD", x"36", x"07", x"FF", x"DD", x"36", x"08", x"FF", -- 0x4E10,
      x"DD", x"36", x"09", x"FF", x"DD", x"36", x"FB", x"01", -- 0x4E18,
      x"21", x"0B", x"00", x"39", x"01", x"04", x"00", x"ED", -- 0x4E20,
      x"B0", x"DD", x"6E", x"FB", x"DD", x"F9", x"DD", x"E1", -- 0x4E28,
      x"C9", x"CD", x"13", x"3F", x"21", x"EF", x"FF", x"39", -- 0x4E30,
      x"F9", x"DD", x"7E", x"06", x"DD", x"77", x"EF", x"DD", -- 0x4E38,
      x"7E", x"07", x"DD", x"77", x"F0", x"E1", x"E5", x"7E", -- 0x4E40,
      x"DD", x"77", x"FC", x"23", x"7E", x"DD", x"77", x"FD", -- 0x4E48,
      x"DD", x"7E", x"04", x"DD", x"77", x"F1", x"DD", x"7E", -- 0x4E50,
      x"05", x"DD", x"77", x"F2", x"DD", x"6E", x"F1", x"DD", -- 0x4E58,
      x"66", x"F2", x"4E", x"23", x"66", x"69", x"11", x"0A", -- 0x4E60,
      x"00", x"19", x"7E", x"DD", x"77", x"F3", x"23", x"7E", -- 0x4E68,
      x"DD", x"77", x"F4", x"AF", x"DD", x"77", x"FE", x"AF", -- 0x4E70,
      x"DD", x"77", x"FF", x"DD", x"6E", x"FC", x"DD", x"66", -- 0x4E78,
      x"FD", x"4E", x"DD", x"34", x"FC", x"20", x"03", x"DD", -- 0x4E80,
      x"34", x"FD", x"DD", x"7E", x"FC", x"DD", x"77", x"F5", -- 0x4E88,
      x"DD", x"7E", x"FD", x"DD", x"77", x"F6", x"79", x"DD", -- 0x4E90,
      x"77", x"F7", x"17", x"9F", x"DD", x"77", x"F8", x"DD", -- 0x4E98,
      x"7E", x"F7", x"DD", x"77", x"F9", x"DD", x"7E", x"F8", -- 0x4EA0,
      x"DD", x"77", x"FA", x"DD", x"7E", x"F9", x"D6", x"20", -- 0x4EA8,
      x"DD", x"7E", x"FA", x"DE", x"00", x"3E", x"00", x"17", -- 0x4EB0,
      x"DD", x"77", x"FB", x"B7", x"20", x"37", x"DD", x"7E", -- 0x4EB8,
      x"F9", x"D6", x"2F", x"DD", x"B6", x"FA", x"28", x"2D", -- 0x4EC0,
      x"DD", x"7E", x"FF", x"D6", x"7F", x"38", x"05", x"2E", -- 0x4EC8,
      x"06", x"C3", x"35", x"52", x"DD", x"6E", x"FF", x"DD", -- 0x4ED0,
      x"34", x"FF", x"DD", x"7E", x"FF", x"DD", x"77", x"FE", -- 0x4ED8,
      x"26", x"00", x"29", x"DD", x"5E", x"F3", x"DD", x"56", -- 0x4EE0,
      x"F4", x"19", x"DD", x"7E", x"F7", x"77", x"23", x"DD", -- 0x4EE8,
      x"7E", x"F8", x"77", x"18", x"86", x"E1", x"E5", x"DD", -- 0x4EF0,
      x"7E", x"F5", x"77", x"23", x"DD", x"7E", x"F6", x"77", -- 0x4EF8,
      x"DD", x"7E", x"FB", x"B7", x"28", x"0A", x"DD", x"36", -- 0x4F00,
      x"FC", x"04", x"AF", x"DD", x"77", x"FD", x"18", x"07", -- 0x4F08,
      x"AF", x"DD", x"77", x"FC", x"DD", x"77", x"FD", x"DD", -- 0x4F10,
      x"7E", x"FC", x"DD", x"77", x"FD", x"DD", x"46", x"FE", -- 0x4F18,
      x"DD", x"70", x"FE", x"AF", x"DD", x"77", x"FF", x"78", -- 0x4F20,
      x"B7", x"28", x"21", x"DD", x"6E", x"FE", x"DD", x"66", -- 0x4F28,
      x"FF", x"2B", x"29", x"DD", x"5E", x"F3", x"DD", x"56", -- 0x4F30,
      x"F4", x"19", x"5E", x"23", x"56", x"7B", x"D6", x"20", -- 0x4F38,
      x"B2", x"28", x"06", x"7B", x"D6", x"2E", x"B2", x"20", -- 0x4F40,
      x"03", x"05", x"18", x"D4", x"DD", x"70", x"FA", x"DD", -- 0x4F48,
      x"6E", x"FE", x"DD", x"66", x"FF", x"29", x"DD", x"5E", -- 0x4F50,
      x"F3", x"DD", x"56", x"F4", x"19", x"AF", x"77", x"23", -- 0x4F58,
      x"77", x"78", x"B7", x"20", x"05", x"2E", x"06", x"C3", -- 0x4F60,
      x"35", x"52", x"AF", x"DD", x"77", x"FF", x"DD", x"7E", -- 0x4F68,
      x"FF", x"DD", x"77", x"FB", x"AF", x"DD", x"77", x"FC", -- 0x4F70,
      x"DD", x"7E", x"FB", x"DD", x"77", x"F8", x"DD", x"7E", -- 0x4F78,
      x"FC", x"DD", x"77", x"F9", x"DD", x"CB", x"F8", x"26", -- 0x4F80,
      x"DD", x"CB", x"F9", x"16", x"DD", x"7E", x"F3", x"DD", -- 0x4F88,
      x"86", x"F8", x"DD", x"77", x"FB", x"DD", x"7E", x"F4", -- 0x4F90,
      x"DD", x"8E", x"F9", x"DD", x"77", x"FC", x"DD", x"6E", -- 0x4F98,
      x"FB", x"DD", x"66", x"FC", x"7E", x"DD", x"77", x"FB", -- 0x4FA0,
      x"23", x"7E", x"DD", x"77", x"FC", x"DD", x"7E", x"FB", -- 0x4FA8,
      x"D6", x"20", x"DD", x"B6", x"FC", x"20", x"05", x"DD", -- 0x4FB0,
      x"34", x"FF", x"18", x"B2", x"DD", x"7E", x"FF", x"DD", -- 0x4FB8,
      x"77", x"FE", x"DD", x"7E", x"FF", x"B7", x"20", x"0A", -- 0x4FC0,
      x"DD", x"7E", x"FB", x"D6", x"2E", x"DD", x"B6", x"FC", -- 0x4FC8,
      x"20", x"08", x"DD", x"7E", x"FD", x"F6", x"03", x"DD", -- 0x4FD0,
      x"77", x"FD", x"DD", x"46", x"FA", x"78", x"B7", x"28", -- 0x4FD8,
      x"18", x"68", x"26", x"00", x"2B", x"29", x"DD", x"5E", -- 0x4FE0,
      x"F3", x"DD", x"56", x"F4", x"19", x"5E", x"23", x"56", -- 0x4FE8,
      x"7B", x"D6", x"2E", x"B2", x"28", x"03", x"05", x"18", -- 0x4FF0,
      x"E4", x"DD", x"70", x"F5", x"DD", x"7E", x"F1", x"C6", -- 0x4FF8,
      x"1C", x"DD", x"77", x"F6", x"DD", x"7E", x"F2", x"CE", -- 0x5000,
      x"00", x"DD", x"77", x"F7", x"DD", x"4E", x"F6", x"DD", -- 0x5008,
      x"46", x"F7", x"21", x"0B", x"00", x"E5", x"2E", x"20", -- 0x5010,
      x"E5", x"C5", x"CD", x"D1", x"00", x"F1", x"F1", x"F1", -- 0x5018,
      x"1E", x"00", x"AF", x"DD", x"77", x"FF", x"DD", x"36", -- 0x5020,
      x"F8", x"08", x"DD", x"6E", x"FE", x"DD", x"34", x"FE", -- 0x5028,
      x"26", x"00", x"29", x"DD", x"4E", x"F3", x"DD", x"46", -- 0x5030,
      x"F4", x"09", x"46", x"23", x"56", x"7B", x"87", x"87", -- 0x5038,
      x"DD", x"77", x"F9", x"7A", x"B0", x"CA", x"B3", x"51", -- 0x5040,
      x"DD", x"70", x"FA", x"DD", x"72", x"FB", x"DD", x"7E", -- 0x5048,
      x"FD", x"F6", x"03", x"4F", x"DD", x"7E", x"FA", x"D6", -- 0x5050,
      x"20", x"DD", x"B6", x"FB", x"28", x"1E", x"DD", x"7E", -- 0x5058,
      x"FE", x"DD", x"96", x"F5", x"3E", x"01", x"28", x"01", -- 0x5060,
      x"AF", x"DD", x"77", x"FC", x"DD", x"7E", x"FA", x"D6", -- 0x5068,
      x"2E", x"DD", x"B6", x"FB", x"20", x"0B", x"DD", x"CB", -- 0x5070,
      x"FC", x"46", x"20", x"05", x"DD", x"71", x"FD", x"18", -- 0x5078,
      x"A9", x"DD", x"7E", x"FF", x"DD", x"96", x"F8", x"30", -- 0x5080,
      x"06", x"DD", x"7E", x"FC", x"B7", x"28", x"33", x"DD", -- 0x5088,
      x"7E", x"F8", x"D6", x"0B", x"20", x"06", x"DD", x"71", -- 0x5090,
      x"FD", x"C3", x"B3", x"51", x"DD", x"CB", x"FC", x"46", -- 0x5098,
      x"20", x"03", x"DD", x"71", x"FD", x"DD", x"7E", x"F5", -- 0x50A0,
      x"DD", x"96", x"FE", x"DA", x"B3", x"51", x"DD", x"7E", -- 0x50A8,
      x"F5", x"DD", x"77", x"FE", x"DD", x"36", x"FF", x"08", -- 0x50B0,
      x"DD", x"36", x"F8", x"0B", x"DD", x"5E", x"F9", x"C3", -- 0x50B8,
      x"2A", x"50", x"DD", x"7E", x"FA", x"D6", x"80", x"DD", -- 0x50C0,
      x"7E", x"FB", x"DE", x"00", x"38", x"1A", x"DD", x"7E", -- 0x50C8,
      x"FD", x"F6", x"02", x"DD", x"77", x"FD", x"CB", x"78", -- 0x50D0,
      x"28", x"0E", x"DD", x"4E", x"FA", x"CB", x"B9", x"06", -- 0x50D8,
      x"00", x"21", x"C6", x"36", x"09", x"46", x"16", x"00", -- 0x50E0,
      x"DD", x"70", x"FB", x"DD", x"72", x"FC", x"DD", x"7E", -- 0x50E8,
      x"FD", x"F6", x"03", x"DD", x"77", x"FA", x"DD", x"7E", -- 0x50F0,
      x"FC", x"D6", x"01", x"38", x"4C", x"DD", x"6E", x"F8", -- 0x50F8,
      x"26", x"00", x"2B", x"DD", x"7E", x"FF", x"DD", x"77", -- 0x5100,
      x"FB", x"AF", x"DD", x"77", x"FC", x"DD", x"7E", x"FB", -- 0x5108,
      x"95", x"DD", x"7E", x"FC", x"9C", x"E2", x"1A", x"51", -- 0x5110,
      x"EE", x"80", x"FA", x"2C", x"51", x"DD", x"7E", x"FA", -- 0x5118,
      x"DD", x"77", x"FD", x"DD", x"7E", x"F8", x"DD", x"77", -- 0x5120,
      x"FF", x"C3", x"2A", x"50", x"DD", x"7E", x"FF", x"DD", -- 0x5128,
      x"34", x"FF", x"DD", x"86", x"F6", x"6F", x"3E", x"00", -- 0x5130,
      x"DD", x"8E", x"F7", x"67", x"DD", x"72", x"FB", x"DD", -- 0x5138,
      x"36", x"FC", x"00", x"DD", x"7E", x"FB", x"77", x"18", -- 0x5140,
      x"56", x"7A", x"B0", x"28", x"14", x"68", x"62", x"C5", -- 0x5148,
      x"D5", x"E5", x"21", x"3A", x"52", x"E5", x"CD", x"E7", -- 0x5150,
      x"58", x"F1", x"F1", x"D1", x"C1", x"7C", x"B5", x"28", -- 0x5158,
      x"0A", x"06", x"5F", x"DD", x"7E", x"FA", x"DD", x"77", -- 0x5160,
      x"FD", x"18", x"34", x"DD", x"7E", x"FB", x"D6", x"41", -- 0x5168,
      x"DD", x"7E", x"FC", x"DE", x"00", x"38", x"0E", x"3E", -- 0x5170,
      x"5A", x"DD", x"BE", x"FB", x"3E", x"00", x"DD", x"9E", -- 0x5178,
      x"FC", x"38", x"02", x"CB", x"CB", x"DD", x"7E", x"FB", -- 0x5180,
      x"D6", x"61", x"DD", x"7E", x"FC", x"DE", x"00", x"38", -- 0x5188,
      x"0E", x"3E", x"7A", x"DD", x"BE", x"FB", x"3E", x"00", -- 0x5190,
      x"DD", x"9E", x"FC", x"38", x"02", x"CB", x"C3", x"DD", -- 0x5198,
      x"7E", x"FF", x"DD", x"34", x"FF", x"DD", x"86", x"F6", -- 0x51A0,
      x"6F", x"3E", x"00", x"DD", x"8E", x"F7", x"67", x"70", -- 0x51A8,
      x"C3", x"2A", x"50", x"DD", x"6E", x"F6", x"DD", x"66", -- 0x51B0,
      x"F7", x"7E", x"D6", x"E5", x"20", x"08", x"DD", x"6E", -- 0x51B8,
      x"F6", x"DD", x"66", x"F7", x"36", x"05", x"DD", x"7E", -- 0x51C0,
      x"F8", x"D6", x"08", x"20", x"03", x"DD", x"5E", x"F9", -- 0x51C8,
      x"DD", x"73", x"FE", x"AF", x"DD", x"77", x"FF", x"DD", -- 0x51D0,
      x"7E", x"FE", x"E6", x"0C", x"4F", x"06", x"00", x"79", -- 0x51D8,
      x"D6", x"0C", x"B0", x"28", x"0E", x"DD", x"7E", x"FE", -- 0x51E0,
      x"E6", x"03", x"4F", x"06", x"00", x"79", x"D6", x"03", -- 0x51E8,
      x"B0", x"20", x"08", x"DD", x"7E", x"FD", x"F6", x"02", -- 0x51F0,
      x"DD", x"77", x"FD", x"DD", x"CB", x"FD", x"4E", x"20", -- 0x51F8,
      x"18", x"CB", x"43", x"28", x"08", x"DD", x"7E", x"FD", -- 0x5200,
      x"F6", x"10", x"DD", x"77", x"FD", x"CB", x"53", x"28", -- 0x5208,
      x"08", x"DD", x"7E", x"FD", x"F6", x"08", x"DD", x"77", -- 0x5210,
      x"FD", x"DD", x"7E", x"F1", x"C6", x"27", x"DD", x"77", -- 0x5218,
      x"FE", x"DD", x"7E", x"F2", x"CE", x"00", x"DD", x"77", -- 0x5220,
      x"FF", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"DD", -- 0x5228,
      x"7E", x"FD", x"77", x"2E", x"00", x"DD", x"F9", x"DD", -- 0x5230,
      x"E1", x"C9", x"2B", x"2C", x"3B", x"3D", x"5B", x"5D", -- 0x5238,
      x"00", x"CD", x"13", x"3F", x"F5", x"F5", x"DD", x"4E", -- 0x5240,
      x"04", x"DD", x"46", x"05", x"59", x"50", x"13", x"13", -- 0x5248,
      x"AF", x"12", x"21", x"24", x"00", x"09", x"36", x"FF", -- 0x5250,
      x"23", x"36", x"FF", x"23", x"36", x"FF", x"23", x"36", -- 0x5258,
      x"FF", x"C5", x"DD", x"6E", x"08", x"DD", x"66", x"09", -- 0x5260,
      x"E5", x"DD", x"6E", x"06", x"DD", x"66", x"07", x"E5", -- 0x5268,
      x"C5", x"CD", x"A2", x"4D", x"F1", x"F1", x"F1", x"7D", -- 0x5270,
      x"C1", x"B7", x"28", x"05", x"2E", x"04", x"C3", x"01", -- 0x5278,
      x"53", x"33", x"33", x"C5", x"DD", x"71", x"FE", x"DD", -- 0x5280,
      x"70", x"FF", x"69", x"60", x"11", x"27", x"02", x"19", -- 0x5288,
      x"56", x"1E", x"00", x"DD", x"6E", x"FE", x"DD", x"66", -- 0x5290,
      x"FF", x"C5", x"01", x"26", x"02", x"09", x"C1", x"6E", -- 0x5298,
      x"26", x"00", x"7B", x"B5", x"5F", x"7A", x"B4", x"57", -- 0x52A0,
      x"7B", x"D6", x"55", x"20", x"05", x"7A", x"D6", x"AA", -- 0x52A8,
      x"28", x"04", x"2E", x"03", x"18", x"4B", x"E1", x"E5", -- 0x52B0,
      x"11", x"28", x"00", x"19", x"7E", x"FE", x"E9", x"28", -- 0x52B8,
      x"08", x"FE", x"EB", x"28", x"04", x"D6", x"E8", x"20", -- 0x52C0,
      x"36", x"21", x"5E", x"00", x"09", x"C5", x"11", x"03", -- 0x52C8,
      x"00", x"D5", x"11", x"06", x"53", x"D5", x"E5", x"CD", -- 0x52D0,
      x"F8", x"5B", x"F1", x"F1", x"F1", x"C1", x"7C", x"B5", -- 0x52D8,
      x"20", x"03", x"6F", x"18", x"1C", x"21", x"7A", x"00", -- 0x52E0,
      x"09", x"01", x"05", x"00", x"C5", x"01", x"0A", x"53", -- 0x52E8,
      x"C5", x"E5", x"CD", x"F8", x"5B", x"F1", x"F1", x"F1", -- 0x52F0,
      x"7C", x"B5", x"20", x"03", x"6F", x"18", x"02", x"2E", -- 0x52F8,
      x"02", x"DD", x"F9", x"DD", x"E1", x"C9", x"46", x"41", -- 0x5300,
      x"54", x"00", x"46", x"41", x"54", x"33", x"32", x"00", -- 0x5308,
      x"F1", x"C1", x"D1", x"D5", x"C5", x"F5", x"AF", x"6F", -- 0x5310,
      x"B0", x"06", x"10", x"20", x"04", x"06", x"08", x"79", -- 0x5318,
      x"29", x"CB", x"11", x"17", x"30", x"01", x"19", x"10", -- 0x5320,
      x"F7", x"C9", x"CD", x"13", x"3F", x"21", x"EE", x"FF", -- 0x5328,
      x"39", x"F9", x"DD", x"36", x"F1", x"04", x"DD", x"4E", -- 0x5330,
      x"04", x"DD", x"46", x"05", x"0A", x"DD", x"77", x"F2", -- 0x5338,
      x"03", x"0A", x"DD", x"77", x"F3", x"0B", x"DD", x"36", -- 0x5340,
      x"F4", x"FF", x"DD", x"36", x"F5", x"FF", x"DD", x"71", -- 0x5348,
      x"F6", x"DD", x"70", x"F7", x"DD", x"7E", x"F2", x"DD", -- 0x5350,
      x"77", x"F8", x"DD", x"7E", x"F3", x"DD", x"77", x"F9", -- 0x5358,
      x"21", x"16", x"00", x"09", x"DD", x"75", x"FA", x"DD", -- 0x5360,
      x"74", x"FB", x"C5", x"DD", x"5E", x"FA", x"DD", x"56", -- 0x5368,
      x"FB", x"21", x"10", x"00", x"39", x"EB", x"01", x"04", -- 0x5370,
      x"00", x"ED", x"B0", x"C1", x"DD", x"7E", x"FF", x"DD", -- 0x5378,
      x"B6", x"FE", x"DD", x"B6", x"FD", x"DD", x"B6", x"FC", -- 0x5380,
      x"CA", x"05", x"55", x"C5", x"DD", x"6E", x"FE", x"DD", -- 0x5388,
      x"66", x"FF", x"E5", x"DD", x"6E", x"FC", x"DD", x"66", -- 0x5390,
      x"FD", x"E5", x"DD", x"6E", x"F2", x"DD", x"66", x"F3", -- 0x5398,
      x"E5", x"CD", x"A2", x"4D", x"F1", x"F1", x"F1", x"C1", -- 0x53A0,
      x"DD", x"75", x"F1", x"7D", x"B7", x"C2", x"05", x"55", -- 0x53A8,
      x"21", x"1A", x"00", x"09", x"DD", x"75", x"FC", x"DD", -- 0x53B0,
      x"74", x"FD", x"7E", x"23", x"66", x"6F", x"7E", x"DD", -- 0x53B8,
      x"77", x"FF", x"B7", x"20", x"07", x"DD", x"36", x"F1", -- 0x53C0,
      x"04", x"C3", x"05", x"55", x"79", x"C6", x"04", x"5F", -- 0x53C8,
      x"78", x"CE", x"00", x"57", x"C5", x"01", x"0B", x"00", -- 0x53D0,
      x"09", x"C1", x"7E", x"E6", x"3F", x"DD", x"77", x"FE", -- 0x53D8,
      x"12", x"DD", x"7E", x"FF", x"D6", x"E5", x"28", x"25", -- 0x53E0,
      x"DD", x"7E", x"FF", x"D6", x"2E", x"28", x"1E", x"DD", -- 0x53E8,
      x"5E", x"FE", x"16", x"00", x"CB", x"AB", x"7B", x"D6", -- 0x53F0,
      x"08", x"B2", x"3E", x"01", x"28", x"01", x"AF", x"5F", -- 0x53F8,
      x"16", x"00", x"DD", x"6E", x"06", x"DD", x"66", x"07", -- 0x5400,
      x"BF", x"ED", x"52", x"28", x"07", x"DD", x"36", x"F4", -- 0x5408,
      x"FF", x"C3", x"F1", x"54", x"21", x"28", x"00", x"09", -- 0x5410,
      x"EB", x"DD", x"7E", x"FE", x"D6", x"0F", x"C2", x"C3", -- 0x5418,
      x"54", x"DD", x"CB", x"FF", x"76", x"28", x"49", x"DD", -- 0x5420,
      x"6E", x"FC", x"DD", x"66", x"FD", x"7E", x"23", x"66", -- 0x5428,
      x"6F", x"C5", x"01", x"0D", x"00", x"09", x"C1", x"7E", -- 0x5430,
      x"DD", x"77", x"F5", x"DD", x"7E", x"FF", x"E6", x"BF", -- 0x5438,
      x"DD", x"77", x"FF", x"DD", x"77", x"F4", x"DD", x"6E", -- 0x5440,
      x"F6", x"DD", x"66", x"F7", x"C5", x"01", x"0E", x"00", -- 0x5448,
      x"09", x"C1", x"7E", x"DD", x"77", x"EE", x"23", x"7E", -- 0x5450,
      x"DD", x"77", x"EF", x"23", x"7E", x"DD", x"77", x"F0", -- 0x5458,
      x"23", x"7E", x"DD", x"77", x"F1", x"C5", x"21", x"02", -- 0x5460,
      x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", x"C1", -- 0x5468,
      x"DD", x"7E", x"F4", x"DD", x"96", x"FF", x"20", x"43", -- 0x5470,
      x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"5E", x"23", -- 0x5478,
      x"56", x"6B", x"62", x"C5", x"01", x"0D", x"00", x"09", -- 0x5480,
      x"C1", x"7E", x"DD", x"77", x"FF", x"DD", x"7E", x"F5", -- 0x5488,
      x"DD", x"96", x"FF", x"20", x"26", x"DD", x"6E", x"F8", -- 0x5490,
      x"DD", x"66", x"F9", x"C5", x"01", x"0A", x"00", x"09", -- 0x5498,
      x"C1", x"7E", x"23", x"66", x"6F", x"C5", x"D5", x"E5", -- 0x54A0,
      x"CD", x"BF", x"57", x"F1", x"F1", x"C1", x"7C", x"B5", -- 0x54A8,
      x"28", x"09", x"DD", x"7E", x"F4", x"3D", x"5F", x"17", -- 0x54B0,
      x"9F", x"18", x"03", x"11", x"FF", x"00", x"DD", x"73", -- 0x54B8,
      x"F4", x"18", x"2E", x"DD", x"7E", x"F4", x"B7", x"20", -- 0x54C0,
      x"17", x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"4E", -- 0x54C8,
      x"23", x"46", x"D5", x"C5", x"CD", x"21", x"55", x"F1", -- 0x54D0,
      x"4D", x"D1", x"DD", x"7E", x"F5", x"91", x"28", x"25", -- 0x54D8,
      x"3E", x"FF", x"12", x"13", x"3E", x"FF", x"12", x"13", -- 0x54E0,
      x"3E", x"FF", x"12", x"13", x"3E", x"FF", x"12", x"18", -- 0x54E8,
      x"14", x"C5", x"21", x"00", x"00", x"E5", x"C5", x"CD", -- 0x54F0,
      x"0B", x"59", x"F1", x"F1", x"C1", x"DD", x"75", x"F1", -- 0x54F8,
      x"7D", x"B7", x"CA", x"6A", x"53", x"DD", x"7E", x"F1", -- 0x5500,
      x"B7", x"28", x"0E", x"DD", x"6E", x"FA", x"DD", x"66", -- 0x5508,
      x"FB", x"AF", x"77", x"23", x"77", x"23", x"77", x"23", -- 0x5510,
      x"77", x"DD", x"6E", x"F1", x"DD", x"F9", x"DD", x"E1", -- 0x5518,
      x"C9", x"CD", x"13", x"3F", x"3B", x"AF", x"DD", x"77", -- 0x5520,
      x"FF", x"01", x"0B", x"00", x"DD", x"6E", x"04", x"DD", -- 0x5528,
      x"66", x"05", x"DD", x"5E", x"FF", x"CB", x"3B", x"DD", -- 0x5530,
      x"7E", x"FF", x"0F", x"E6", x"80", x"83", x"5E", x"23", -- 0x5538,
      x"83", x"DD", x"77", x"FF", x"59", x"50", x"1B", x"4B", -- 0x5540,
      x"7A", x"47", x"B3", x"20", x"E5", x"DD", x"6E", x"FF", -- 0x5548,
      x"33", x"DD", x"E1", x"C9", x"CD", x"13", x"3F", x"21", -- 0x5550,
      x"E5", x"FF", x"39", x"F9", x"DD", x"7E", x"04", x"DD", -- 0x5558,
      x"77", x"FE", x"DD", x"7E", x"05", x"DD", x"77", x"FF", -- 0x5560,
      x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"7E", x"DD", -- 0x5568,
      x"77", x"E9", x"23", x"7E", x"DD", x"77", x"EA", x"21", -- 0x5570,
      x"00", x"00", x"E5", x"21", x"00", x"00", x"E5", x"DD", -- 0x5578,
      x"6E", x"FE", x"DD", x"66", x"FF", x"E5", x"CD", x"B6", -- 0x5580,
      x"46", x"F1", x"F1", x"F1", x"DD", x"75", x"FD", x"7D", -- 0x5588,
      x"B7", x"28", x"06", x"DD", x"6E", x"FD", x"C3", x"BA", -- 0x5590,
      x"57", x"DD", x"36", x"EB", x"FF", x"DD", x"36", x"EC", -- 0x5598,
      x"FF", x"DD", x"7E", x"FE", x"DD", x"77", x"ED", x"DD", -- 0x55A0,
      x"7E", x"FF", x"DD", x"77", x"EE", x"DD", x"7E", x"FE", -- 0x55A8,
      x"C6", x"28", x"DD", x"77", x"EF", x"DD", x"7E", x"FF", -- 0x55B0,
      x"CE", x"00", x"DD", x"77", x"F0", x"DD", x"6E", x"EF", -- 0x55B8,
      x"DD", x"66", x"F0", x"36", x"FF", x"23", x"36", x"FF", -- 0x55C0,
      x"23", x"36", x"FF", x"23", x"36", x"FF", x"DD", x"7E", -- 0x55C8,
      x"FE", x"DD", x"77", x"F1", x"DD", x"7E", x"FF", x"DD", -- 0x55D0,
      x"77", x"F2", x"DD", x"7E", x"E9", x"DD", x"77", x"F3", -- 0x55D8,
      x"DD", x"7E", x"EA", x"DD", x"77", x"F4", x"DD", x"7E", -- 0x55E0,
      x"FE", x"C6", x"1C", x"DD", x"77", x"F5", x"DD", x"7E", -- 0x55E8,
      x"FF", x"CE", x"00", x"DD", x"77", x"F6", x"DD", x"7E", -- 0x55F0,
      x"FE", x"C6", x"27", x"DD", x"77", x"F7", x"DD", x"7E", -- 0x55F8,
      x"FF", x"CE", x"00", x"DD", x"77", x"F8", x"DD", x"7E", -- 0x5600,
      x"F7", x"DD", x"77", x"F9", x"DD", x"7E", x"F8", x"DD", -- 0x5608,
      x"77", x"FA", x"DD", x"7E", x"FE", x"DD", x"77", x"FB", -- 0x5610,
      x"DD", x"7E", x"FF", x"DD", x"77", x"FC", x"DD", x"6E", -- 0x5618,
      x"FB", x"DD", x"66", x"FC", x"11", x"16", x"00", x"19", -- 0x5620,
      x"4E", x"23", x"46", x"23", x"5E", x"23", x"56", x"D5", -- 0x5628,
      x"C5", x"DD", x"6E", x"E9", x"DD", x"66", x"EA", x"E5", -- 0x5630,
      x"CD", x"A2", x"4D", x"F1", x"F1", x"F1", x"DD", x"75", -- 0x5638,
      x"FD", x"7D", x"B7", x"C2", x"B7", x"57", x"DD", x"7E", -- 0x5640,
      x"ED", x"C6", x"1A", x"4F", x"DD", x"7E", x"EE", x"CE", -- 0x5648,
      x"00", x"47", x"69", x"60", x"7E", x"23", x"66", x"6F", -- 0x5650,
      x"5E", x"7B", x"B7", x"20", x"07", x"DD", x"36", x"FD", -- 0x5658,
      x"04", x"C3", x"B7", x"57", x"DD", x"7E", x"ED", x"C6", -- 0x5660,
      x"04", x"DD", x"77", x"FE", x"DD", x"7E", x"EE", x"CE", -- 0x5668,
      x"00", x"DD", x"77", x"FF", x"C5", x"01", x"0B", x"00", -- 0x5670,
      x"09", x"C1", x"7E", x"E6", x"3F", x"57", x"DD", x"6E", -- 0x5678,
      x"FE", x"DD", x"66", x"FF", x"77", x"7B", x"D6", x"E5", -- 0x5680,
      x"28", x"10", x"7A", x"D6", x"0F", x"3E", x"01", x"28", -- 0x5688,
      x"01", x"AF", x"CB", x"5A", x"28", x"1C", x"CB", x"47", -- 0x5690,
      x"20", x"18", x"DD", x"36", x"EC", x"FF", x"DD", x"6E", -- 0x5698,
      x"EF", x"DD", x"66", x"F0", x"36", x"FF", x"23", x"36", -- 0x56A0,
      x"FF", x"23", x"36", x"FF", x"23", x"36", x"FF", x"C3", -- 0x56A8,
      x"9F", x"57", x"B7", x"CA", x"4C", x"57", x"DD", x"6E", -- 0x56B0,
      x"F9", x"DD", x"66", x"FA", x"CB", x"76", x"C2", x"9F", -- 0x56B8,
      x"57", x"CB", x"73", x"28", x"47", x"69", x"60", x"56", -- 0x56C0,
      x"23", x"66", x"6A", x"C5", x"01", x"0D", x"00", x"09", -- 0x56C8,
      x"C1", x"7E", x"DD", x"77", x"EB", x"CB", x"B3", x"DD", -- 0x56D0,
      x"73", x"EC", x"DD", x"6E", x"F1", x"DD", x"66", x"F2", -- 0x56D8,
      x"C5", x"01", x"0E", x"00", x"09", x"C1", x"7E", x"DD", -- 0x56E0,
      x"77", x"E5", x"23", x"7E", x"DD", x"77", x"E6", x"23", -- 0x56E8,
      x"7E", x"DD", x"77", x"E7", x"23", x"7E", x"DD", x"77", -- 0x56F0,
      x"E8", x"D5", x"C5", x"DD", x"5E", x"EF", x"DD", x"56", -- 0x56F8,
      x"F0", x"21", x"04", x"00", x"39", x"01", x"04", x"00", -- 0x5700,
      x"ED", x"B0", x"C1", x"D1", x"DD", x"7E", x"EC", x"93", -- 0x5708,
      x"20", x"32", x"69", x"60", x"5E", x"23", x"56", x"6B", -- 0x5710,
      x"62", x"01", x"0D", x"00", x"09", x"DD", x"7E", x"EB", -- 0x5718,
      x"96", x"20", x"21", x"DD", x"6E", x"F3", x"DD", x"66", -- 0x5720,
      x"F4", x"01", x"0A", x"00", x"09", x"4E", x"23", x"46", -- 0x5728,
      x"D5", x"C5", x"CD", x"47", x"5C", x"F1", x"F1", x"7C", -- 0x5730,
      x"B5", x"28", x"09", x"DD", x"7E", x"EC", x"3D", x"4F", -- 0x5738,
      x"17", x"9F", x"18", x"03", x"01", x"FF", x"00", x"DD", -- 0x5740,
      x"71", x"EC", x"18", x"53", x"DD", x"7E", x"EC", x"B7", -- 0x5748,
      x"20", x"13", x"69", x"60", x"5E", x"23", x"56", x"C5", -- 0x5750,
      x"D5", x"CD", x"21", x"55", x"F1", x"5D", x"C1", x"DD", -- 0x5758,
      x"7E", x"EB", x"93", x"28", x"52", x"DD", x"6E", x"F7", -- 0x5760,
      x"DD", x"66", x"F8", x"7E", x"0F", x"38", x"1B", x"DD", -- 0x5768,
      x"5E", x"F5", x"DD", x"56", x"F6", x"69", x"60", x"4E", -- 0x5770,
      x"23", x"46", x"21", x"0B", x"00", x"E5", x"D5", x"C5", -- 0x5778,
      x"CD", x"F8", x"5B", x"F1", x"F1", x"F1", x"7C", x"B5", -- 0x5780,
      x"28", x"2D", x"DD", x"36", x"EC", x"FF", x"DD", x"6E", -- 0x5788,
      x"EF", x"DD", x"66", x"F0", x"36", x"FF", x"23", x"36", -- 0x5790,
      x"FF", x"23", x"36", x"FF", x"23", x"36", x"FF", x"21", -- 0x5798,
      x"00", x"00", x"E5", x"DD", x"6E", x"ED", x"DD", x"66", -- 0x57A0,
      x"EE", x"E5", x"CD", x"0B", x"59", x"F1", x"F1", x"DD", -- 0x57A8,
      x"75", x"FD", x"7D", x"B7", x"CA", x"1E", x"56", x"DD", -- 0x57B0,
      x"6E", x"FD", x"DD", x"F9", x"DD", x"E1", x"C9", x"CD", -- 0x57B8,
      x"13", x"3F", x"21", x"F6", x"FF", x"39", x"F9", x"DD", -- 0x57C0,
      x"7E", x"06", x"C6", x"1A", x"5F", x"DD", x"7E", x"07", -- 0x57C8,
      x"CE", x"00", x"57", x"6B", x"62", x"23", x"46", x"0E", -- 0x57D0,
      x"00", x"1A", x"5F", x"16", x"00", x"79", x"B3", x"4F", -- 0x57D8,
      x"78", x"B2", x"B1", x"28", x"06", x"21", x"00", x"00", -- 0x57E0,
      x"C3", x"E2", x"58", x"DD", x"7E", x"06", x"DD", x"77", -- 0x57E8,
      x"F6", x"DD", x"7E", x"07", x"DD", x"77", x"F7", x"E1", -- 0x57F0,
      x"E5", x"4E", x"06", x"00", x"CB", x"B1", x"0B", x"69", -- 0x57F8,
      x"60", x"29", x"09", x"29", x"29", x"09", x"DD", x"75", -- 0x5800,
      x"F8", x"DD", x"74", x"F9", x"DD", x"36", x"FA", x"01", -- 0x5808,
      x"AF", x"DD", x"77", x"FB", x"DD", x"7E", x"F8", x"DD", -- 0x5810,
      x"77", x"FE", x"DD", x"7E", x"F9", x"DD", x"77", x"FF", -- 0x5818,
      x"01", x"00", x"00", x"79", x"D6", x"0D", x"78", x"DE", -- 0x5820,
      x"00", x"D2", x"B5", x"58", x"21", x"B9", x"36", x"09", -- 0x5828,
      x"7E", x"DD", x"86", x"F6", x"5F", x"3E", x"00", x"DD", -- 0x5830,
      x"8E", x"F7", x"57", x"6B", x"62", x"23", x"6E", x"DD", -- 0x5838,
      x"75", x"FD", x"DD", x"36", x"FC", x"00", x"1A", x"5F", -- 0x5840,
      x"16", x"00", x"DD", x"7E", x"FC", x"B3", x"5F", x"DD", -- 0x5848,
      x"7E", x"FD", x"B2", x"57", x"DD", x"7E", x"FB", x"DD", -- 0x5850,
      x"B6", x"FA", x"28", x"4B", x"DD", x"7E", x"FE", x"D6", -- 0x5858,
      x"7F", x"DD", x"7E", x"FF", x"DE", x"00", x"38", x"05", -- 0x5860,
      x"21", x"00", x"00", x"18", x"75", x"DD", x"6E", x"FE", -- 0x5868,
      x"DD", x"66", x"FF", x"DD", x"34", x"FE", x"20", x"03", -- 0x5870,
      x"DD", x"34", x"FF", x"DD", x"7E", x"FE", x"DD", x"77", -- 0x5878,
      x"F8", x"DD", x"7E", x"FF", x"DD", x"77", x"F9", x"29", -- 0x5880,
      x"DD", x"75", x"FC", x"DD", x"74", x"FD", x"DD", x"7E", -- 0x5888,
      x"04", x"DD", x"86", x"FC", x"6F", x"DD", x"7E", x"05", -- 0x5890,
      x"DD", x"8E", x"FD", x"67", x"DD", x"73", x"FA", x"DD", -- 0x5898,
      x"72", x"FB", x"73", x"23", x"72", x"18", x"0A", x"7B", -- 0x58A0,
      x"A2", x"3C", x"28", x"05", x"21", x"00", x"00", x"18", -- 0x58A8,
      x"31", x"03", x"C3", x"23", x"58", x"E1", x"E5", x"CB", -- 0x58B0,
      x"76", x"28", x"24", x"DD", x"7E", x"F8", x"D6", x"7F", -- 0x58B8,
      x"DD", x"7E", x"F9", x"DE", x"00", x"38", x"05", x"21", -- 0x58C0,
      x"00", x"00", x"18", x"16", x"D1", x"C1", x"C5", x"D5", -- 0x58C8,
      x"CB", x"21", x"CB", x"10", x"DD", x"6E", x"04", x"DD", -- 0x58D0,
      x"66", x"05", x"09", x"AF", x"77", x"23", x"77", x"21", -- 0x58D8,
      x"01", x"00", x"DD", x"F9", x"DD", x"E1", x"C9", x"D1", -- 0x58E0,
      x"C1", x"C5", x"D5", x"0A", x"F5", x"5F", x"17", x"9F", -- 0x58E8,
      x"57", x"F1", x"B7", x"28", x"14", x"FD", x"21", x"04", -- 0x58F0,
      x"00", x"FD", x"39", x"FD", x"6E", x"00", x"FD", x"66", -- 0x58F8,
      x"01", x"BF", x"ED", x"52", x"28", x"03", x"03", x"18", -- 0x5900,
      x"E2", x"EB", x"C9", x"CD", x"13", x"3F", x"21", x"E6", -- 0x5908,
      x"FF", x"39", x"F9", x"DD", x"7E", x"04", x"DD", x"77", -- 0x5910,
      x"E6", x"DD", x"7E", x"05", x"DD", x"77", x"E7", x"E1", -- 0x5918,
      x"E5", x"7E", x"DD", x"77", x"E8", x"23", x"7E", x"DD", -- 0x5920,
      x"77", x"E9", x"DD", x"7E", x"E6", x"C6", x"0E", x"DD", -- 0x5928,
      x"77", x"EA", x"DD", x"7E", x"E7", x"CE", x"00", x"DD", -- 0x5930,
      x"77", x"EB", x"DD", x"6E", x"EA", x"DD", x"66", x"EB", -- 0x5938,
      x"4E", x"23", x"46", x"23", x"5E", x"23", x"56", x"79", -- 0x5940,
      x"C6", x"20", x"DD", x"77", x"EC", x"78", x"CE", x"00", -- 0x5948,
      x"DD", x"77", x"ED", x"7B", x"CE", x"00", x"DD", x"77", -- 0x5950,
      x"EE", x"7A", x"CE", x"00", x"DD", x"77", x"EF", x"DD", -- 0x5958,
      x"7E", x"E6", x"C6", x"16", x"DD", x"77", x"F0", x"DD", -- 0x5960,
      x"7E", x"E7", x"CE", x"00", x"DD", x"77", x"F1", x"DD", -- 0x5968,
      x"7E", x"EE", x"D6", x"20", x"DD", x"7E", x"EF", x"DE", -- 0x5970,
      x"00", x"38", x"0E", x"DD", x"6E", x"F0", x"DD", x"66", -- 0x5978,
      x"F1", x"AF", x"77", x"23", x"77", x"23", x"77", x"23", -- 0x5980,
      x"77", x"DD", x"5E", x"F0", x"DD", x"56", x"F1", x"21", -- 0x5988,
      x"16", x"00", x"39", x"EB", x"01", x"04", x"00", x"ED", -- 0x5990,
      x"B0", x"DD", x"7E", x"FF", x"DD", x"B6", x"FE", x"DD", -- 0x5998,
      x"B6", x"FD", x"DD", x"B6", x"FC", x"20", x"05", x"2E", -- 0x59A0,
      x"04", x"C3", x"F3", x"5B", x"DD", x"7E", x"EC", x"DD", -- 0x59A8,
      x"77", x"F2", x"DD", x"7E", x"ED", x"E6", x"01", x"DD", -- 0x59B0,
      x"77", x"F3", x"DD", x"36", x"F4", x"00", x"DD", x"36", -- 0x59B8,
      x"F5", x"00", x"3E", x"00", x"DD", x"B6", x"F4", x"DD", -- 0x59C0,
      x"B6", x"F3", x"DD", x"B6", x"F2", x"C2", x"A1", x"5B", -- 0x59C8,
      x"DD", x"7E", x"FC", x"C6", x"01", x"4F", x"DD", x"7E", -- 0x59D0,
      x"FD", x"CE", x"00", x"47", x"DD", x"7E", x"FE", x"CE", -- 0x59D8,
      x"00", x"5F", x"DD", x"7E", x"FF", x"CE", x"00", x"57", -- 0x59E0,
      x"DD", x"6E", x"F0", x"DD", x"66", x"F1", x"71", x"23", -- 0x59E8,
      x"70", x"23", x"73", x"23", x"72", x"DD", x"7E", x"E6", -- 0x59F0,
      x"C6", x"12", x"DD", x"77", x"F6", x"DD", x"7E", x"E7", -- 0x59F8,
      x"CE", x"00", x"DD", x"77", x"F7", x"DD", x"5E", x"F6", -- 0x5A00,
      x"DD", x"56", x"F7", x"21", x"12", x"00", x"39", x"EB", -- 0x5A08,
      x"01", x"04", x"00", x"ED", x"B0", x"DD", x"7E", x"FB", -- 0x5A10,
      x"DD", x"B6", x"FA", x"DD", x"B6", x"F9", x"DD", x"B6", -- 0x5A18,
      x"F8", x"20", x"5B", x"DD", x"4E", x"EC", x"DD", x"46", -- 0x5A20,
      x"ED", x"DD", x"5E", x"EE", x"DD", x"56", x"EF", x"3E", -- 0x5A28,
      x"05", x"CB", x"3A", x"CB", x"1B", x"CB", x"18", x"CB", -- 0x5A30,
      x"19", x"3D", x"20", x"F5", x"DD", x"6E", x"E8", x"DD", -- 0x5A38,
      x"66", x"E9", x"C5", x"01", x"06", x"00", x"09", x"C1", -- 0x5A40,
      x"7E", x"23", x"66", x"DD", x"77", x"FC", x"DD", x"74", -- 0x5A48,
      x"FD", x"AF", x"DD", x"77", x"FE", x"DD", x"77", x"FF", -- 0x5A50,
      x"79", x"DD", x"96", x"FC", x"78", x"DD", x"9E", x"FD", -- 0x5A58,
      x"7B", x"DD", x"9E", x"FE", x"7A", x"DD", x"9E", x"FF", -- 0x5A60,
      x"DA", x"A1", x"5B", x"DD", x"6E", x"F0", x"DD", x"66", -- 0x5A68,
      x"F1", x"AF", x"77", x"23", x"77", x"23", x"77", x"23", -- 0x5A70,
      x"77", x"2E", x"04", x"C3", x"F3", x"5B", x"DD", x"4E", -- 0x5A78,
      x"ED", x"DD", x"46", x"EE", x"DD", x"5E", x"EF", x"16", -- 0x5A80,
      x"00", x"CB", x"3B", x"CB", x"18", x"CB", x"19", x"DD", -- 0x5A88,
      x"6E", x"E8", x"DD", x"66", x"E9", x"C5", x"01", x"09", -- 0x5A90,
      x"00", x"09", x"C1", x"7E", x"2B", x"6E", x"67", x"2B", -- 0x5A98,
      x"DD", x"75", x"FC", x"DD", x"74", x"FD", x"AF", x"DD", -- 0x5AA0,
      x"77", x"FE", x"DD", x"77", x"FF", x"79", x"DD", x"A6", -- 0x5AA8,
      x"FC", x"F5", x"78", x"DD", x"A6", x"FD", x"4F", x"7B", -- 0x5AB0,
      x"DD", x"A6", x"FE", x"6F", x"7A", x"DD", x"A6", x"FF", -- 0x5AB8,
      x"67", x"F1", x"B4", x"B5", x"B1", x"C2", x"A1", x"5B", -- 0x5AC0,
      x"DD", x"6E", x"FA", x"DD", x"66", x"FB", x"E5", x"DD", -- 0x5AC8,
      x"6E", x"F8", x"DD", x"66", x"F9", x"E5", x"DD", x"6E", -- 0x5AD0,
      x"E6", x"DD", x"66", x"E7", x"E5", x"CD", x"C1", x"44", -- 0x5AD8,
      x"F1", x"F1", x"F1", x"DD", x"75", x"FC", x"DD", x"74", -- 0x5AE0,
      x"FD", x"DD", x"73", x"FE", x"DD", x"72", x"FF", x"3E", -- 0x5AE8,
      x"01", x"DD", x"BE", x"FC", x"3E", x"00", x"DD", x"9E", -- 0x5AF0,
      x"FD", x"3E", x"00", x"DD", x"9E", x"FE", x"3E", x"00", -- 0x5AF8,
      x"DD", x"9E", x"FF", x"38", x"05", x"2E", x"02", x"C3", -- 0x5B00,
      x"F3", x"5B", x"DD", x"7E", x"FC", x"DD", x"A6", x"FD", -- 0x5B08,
      x"DD", x"A6", x"FE", x"DD", x"A6", x"FF", x"3C", x"20", -- 0x5B10,
      x"05", x"2E", x"01", x"C3", x"F3", x"5B", x"C1", x"E1", -- 0x5B18,
      x"E5", x"C5", x"11", x"0C", x"00", x"19", x"4E", x"23", -- 0x5B20,
      x"46", x"23", x"5E", x"23", x"56", x"DD", x"7E", x"FC", -- 0x5B28,
      x"91", x"DD", x"7E", x"FD", x"98", x"DD", x"7E", x"FE", -- 0x5B30,
      x"9B", x"DD", x"7E", x"FF", x"9A", x"38", x"29", x"DD", -- 0x5B38,
      x"7E", x"07", x"DD", x"B6", x"06", x"20", x"0E", x"DD", -- 0x5B40,
      x"6E", x"F0", x"DD", x"66", x"F1", x"AF", x"77", x"23", -- 0x5B48,
      x"77", x"23", x"77", x"23", x"77", x"DD", x"6E", x"F0", -- 0x5B50,
      x"DD", x"66", x"F1", x"AF", x"77", x"23", x"77", x"23", -- 0x5B58,
      x"77", x"23", x"77", x"2E", x"04", x"C3", x"F3", x"5B", -- 0x5B60,
      x"DD", x"5E", x"F6", x"DD", x"56", x"F7", x"21", x"16", -- 0x5B68,
      x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", x"DD", -- 0x5B70,
      x"6E", x"FE", x"DD", x"66", x"FF", x"E5", x"DD", x"6E", -- 0x5B78,
      x"FC", x"DD", x"66", x"FD", x"E5", x"DD", x"6E", x"E8", -- 0x5B80,
      x"DD", x"66", x"E9", x"E5", x"CD", x"68", x"37", x"F1", -- 0x5B88,
      x"F1", x"F1", x"4D", x"44", x"DD", x"6E", x"F0", x"DD", -- 0x5B90,
      x"66", x"F1", x"71", x"23", x"70", x"23", x"73", x"23", -- 0x5B98,
      x"72", x"DD", x"5E", x"EA", x"DD", x"56", x"EB", x"21", -- 0x5BA0,
      x"06", x"00", x"39", x"01", x"04", x"00", x"ED", x"B0", -- 0x5BA8,
      x"DD", x"7E", x"E6", x"C6", x"1A", x"DD", x"77", x"FE", -- 0x5BB0,
      x"DD", x"7E", x"E7", x"CE", x"00", x"DD", x"77", x"FF", -- 0x5BB8,
      x"DD", x"7E", x"E8", x"C6", x"28", x"DD", x"77", x"FC", -- 0x5BC0,
      x"DD", x"7E", x"E9", x"CE", x"00", x"DD", x"77", x"FD", -- 0x5BC8,
      x"DD", x"7E", x"FC", x"DD", x"86", x"F2", x"DD", x"77", -- 0x5BD0,
      x"FA", x"DD", x"7E", x"FD", x"DD", x"8E", x"F3", x"DD", -- 0x5BD8,
      x"77", x"FB", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", -- 0x5BE0,
      x"DD", x"7E", x"FA", x"77", x"23", x"DD", x"7E", x"FB", -- 0x5BE8,
      x"77", x"2E", x"00", x"DD", x"F9", x"DD", x"E1", x"C9", -- 0x5BF0,
      x"CD", x"13", x"3F", x"F5", x"F5", x"DD", x"4E", x"04", -- 0x5BF8,
      x"DD", x"46", x"05", x"DD", x"7E", x"06", x"DD", x"77", -- 0x5C00,
      x"FE", x"DD", x"7E", x"07", x"DD", x"77", x"FF", x"DD", -- 0x5C08,
      x"5E", x"08", x"DD", x"56", x"09", x"0A", x"03", x"DD", -- 0x5C10,
      x"77", x"FC", x"AF", x"DD", x"77", x"FD", x"DD", x"6E", -- 0x5C18,
      x"FE", x"DD", x"66", x"FF", x"6E", x"DD", x"34", x"FE", -- 0x5C20,
      x"20", x"03", x"DD", x"34", x"FF", x"26", x"00", x"DD", -- 0x5C28,
      x"7E", x"FC", x"95", x"6F", x"DD", x"7E", x"FD", x"9C", -- 0x5C30,
      x"67", x"1B", x"7A", x"B3", x"28", x"04", x"7C", x"B5", -- 0x5C38,
      x"28", x"D3", x"DD", x"F9", x"DD", x"E1", x"C9", x"CD", -- 0x5C40,
      x"13", x"3F", x"21", x"F5", x"FF", x"39", x"F9", x"DD", -- 0x5C48,
      x"7E", x"06", x"C6", x"1A", x"5F", x"DD", x"7E", x"07", -- 0x5C50,
      x"CE", x"00", x"57", x"6B", x"62", x"23", x"46", x"0E", -- 0x5C58,
      x"00", x"1A", x"5F", x"16", x"00", x"79", x"B3", x"4F", -- 0x5C60,
      x"78", x"B2", x"B1", x"28", x"06", x"21", x"00", x"00", -- 0x5C68,
      x"C3", x"84", x"5D", x"DD", x"4E", x"06", x"DD", x"46", -- 0x5C70,
      x"07", x"0A", x"DD", x"77", x"F5", x"E6", x"3F", x"5F", -- 0x5C78,
      x"16", x"00", x"1B", x"6B", x"62", x"29", x"19", x"29", -- 0x5C80,
      x"29", x"19", x"DD", x"75", x"F6", x"DD", x"74", x"F7", -- 0x5C88,
      x"11", x"01", x"00", x"DD", x"7E", x"F6", x"DD", x"77", -- 0x5C90,
      x"FC", x"DD", x"7E", x"F7", x"DD", x"77", x"FD", x"AF", -- 0x5C98,
      x"DD", x"77", x"FE", x"DD", x"77", x"FF", x"DD", x"7E", -- 0x5CA0,
      x"FE", x"D6", x"0D", x"DD", x"7E", x"FF", x"DE", x"00", -- 0x5CA8,
      x"D2", x"5B", x"5D", x"3E", x"B9", x"DD", x"86", x"FE", -- 0x5CB0,
      x"6F", x"3E", x"36", x"DD", x"8E", x"FF", x"67", x"7E", -- 0x5CB8,
      x"81", x"DD", x"77", x"F8", x"3E", x"00", x"88", x"DD", -- 0x5CC0,
      x"77", x"F9", x"DD", x"6E", x"F8", x"DD", x"66", x"F9", -- 0x5CC8,
      x"23", x"6E", x"DD", x"75", x"FB", x"DD", x"36", x"FA", -- 0x5CD0,
      x"00", x"DD", x"6E", x"F8", x"DD", x"66", x"F9", x"6E", -- 0x5CD8,
      x"26", x"00", x"7D", x"DD", x"B6", x"FA", x"6F", x"7C", -- 0x5CE0,
      x"DD", x"B6", x"FB", x"67", x"DD", x"75", x"FA", x"DD", -- 0x5CE8,
      x"74", x"FB", x"7A", x"B3", x"28", x"4A", x"DD", x"7E", -- 0x5CF0,
      x"FC", x"D6", x"7F", x"DD", x"7E", x"FD", x"DE", x"00", -- 0x5CF8,
      x"30", x"31", x"DD", x"6E", x"FC", x"DD", x"66", x"FD", -- 0x5D00,
      x"DD", x"34", x"FC", x"20", x"03", x"DD", x"34", x"FD", -- 0x5D08,
      x"DD", x"7E", x"FC", x"DD", x"77", x"F6", x"DD", x"7E", -- 0x5D10,
      x"FD", x"DD", x"77", x"F7", x"29", x"EB", x"DD", x"6E", -- 0x5D18,
      x"04", x"DD", x"66", x"05", x"19", x"5E", x"23", x"56", -- 0x5D20,
      x"DD", x"6E", x"FA", x"DD", x"66", x"FB", x"BF", x"ED", -- 0x5D28,
      x"52", x"28", x"05", x"21", x"00", x"00", x"18", x"4C", -- 0x5D30,
      x"DD", x"5E", x"FA", x"DD", x"56", x"FB", x"18", x"0F", -- 0x5D38,
      x"DD", x"7E", x"FA", x"DD", x"66", x"FB", x"A4", x"3C", -- 0x5D40,
      x"28", x"05", x"21", x"00", x"00", x"18", x"35", x"DD", -- 0x5D48,
      x"34", x"FE", x"C2", x"A6", x"5C", x"DD", x"34", x"FF", -- 0x5D50,
      x"C3", x"A6", x"5C", x"DD", x"CB", x"F5", x"76", x"28", -- 0x5D58,
      x"20", x"7A", x"B3", x"28", x"1C", x"DD", x"4E", x"F6", -- 0x5D60,
      x"DD", x"46", x"F7", x"CB", x"21", x"CB", x"10", x"DD", -- 0x5D68,
      x"6E", x"04", x"DD", x"66", x"05", x"09", x"7E", x"23", -- 0x5D70,
      x"4E", x"B1", x"28", x"05", x"21", x"00", x"00", x"18", -- 0x5D78,
      x"03", x"21", x"01", x"00", x"DD", x"F9", x"DD", x"E1", -- 0x5D80,
      x"C9", x"DD", x"E5", x"DD", x"21", x"00", x"00", x"DD", -- 0x5D88,
      x"39", x"21", x"F8", x"FF", x"39", x"F9", x"21", x"0C", -- 0x5D90,
      x"00", x"39", x"EB", x"4B", x"42", x"03", x"03", x"DD", -- 0x5D98,
      x"71", x"FE", x"DD", x"70", x"FF", x"6B", x"62", x"23", -- 0x5DA0,
      x"23", x"4E", x"23", x"46", x"21", x"10", x"00", x"39", -- 0x5DA8,
      x"E3", x"E1", x"E5", x"7E", x"23", x"66", x"6F", x"D5", -- 0x5DB0,
      x"E5", x"C5", x"CD", x"10", x"53", x"F1", x"F1", x"4D", -- 0x5DB8,
      x"44", x"D1", x"DD", x"6E", x"FE", x"DD", x"66", x"FF", -- 0x5DC0,
      x"71", x"23", x"70", x"4B", x"42", x"03", x"03", x"DD", -- 0x5DC8,
      x"71", x"FC", x"DD", x"70", x"FD", x"6B", x"62", x"23", -- 0x5DD0,
      x"23", x"7E", x"DD", x"77", x"FE", x"23", x"7E", x"DD", -- 0x5DD8,
      x"77", x"FF", x"E1", x"E5", x"23", x"23", x"4E", x"23", -- 0x5DE0,
      x"46", x"6B", x"62", x"7E", x"23", x"66", x"6F", x"D5", -- 0x5DE8,
      x"E5", x"C5", x"CD", x"10", x"53", x"F1", x"F1", x"D1", -- 0x5DF0,
      x"DD", x"7E", x"FE", x"85", x"4F", x"DD", x"7E", x"FF", -- 0x5DF8,
      x"8C", x"47", x"DD", x"6E", x"FC", x"DD", x"66", x"FD", -- 0x5E00,
      x"71", x"23", x"70", x"4B", x"42", x"03", x"03", x"DD", -- 0x5E08,
      x"71", x"FD", x"DD", x"70", x"FE", x"6B", x"62", x"23", -- 0x5E10,
      x"23", x"4E", x"23", x"46", x"6B", x"62", x"23", x"7E", -- 0x5E18,
      x"DD", x"77", x"FF", x"E1", x"E5", x"23", x"66", x"D5", -- 0x5E20,
      x"C5", x"DD", x"5E", x"FF", x"2E", x"00", x"55", x"06", -- 0x5E28,
      x"08", x"29", x"30", x"01", x"19", x"10", x"FA", x"C1", -- 0x5E30,
      x"D1", x"09", x"4D", x"44", x"DD", x"6E", x"FD", x"DD", -- 0x5E38,
      x"66", x"FE", x"71", x"23", x"70", x"E1", x"E5", x"4E", -- 0x5E40,
      x"6B", x"62", x"23", x"66", x"D5", x"59", x"2E", x"00", -- 0x5E48,
      x"55", x"06", x"08", x"29", x"30", x"01", x"19", x"10", -- 0x5E50,
      x"FA", x"D1", x"DD", x"75", x"FA", x"DD", x"74", x"FB", -- 0x5E58,
      x"C1", x"C5", x"03", x"DD", x"71", x"FE", x"DD", x"70", -- 0x5E60,
      x"FF", x"6B", x"62", x"4E", x"E1", x"E5", x"23", x"66", -- 0x5E68,
      x"D5", x"59", x"2E", x"00", x"55", x"06", x"08", x"29", -- 0x5E70,
      x"30", x"01", x"19", x"10", x"FA", x"D1", x"4D", x"44", -- 0x5E78,
      x"DD", x"6E", x"FE", x"DD", x"66", x"FF", x"71", x"23", -- 0x5E80,
      x"70", x"C1", x"C5", x"03", x"03", x"03", x"DD", x"71", -- 0x5E88,
      x"FC", x"DD", x"70", x"FD", x"C1", x"C5", x"03", x"DD", -- 0x5E90,
      x"71", x"FE", x"DD", x"70", x"FF", x"E1", x"E5", x"23", -- 0x5E98,
      x"4E", x"23", x"46", x"79", x"DD", x"86", x"FA", x"4F", -- 0x5EA0,
      x"78", x"DD", x"8E", x"FB", x"47", x"DD", x"6E", x"FE", -- 0x5EA8,
      x"DD", x"66", x"FF", x"71", x"23", x"70", x"79", x"DD", -- 0x5EB0,
      x"96", x"FA", x"78", x"DD", x"9E", x"FB", x"3E", x"00", -- 0x5EB8,
      x"17", x"DD", x"6E", x"FC", x"DD", x"66", x"FD", x"77", -- 0x5EC0,
      x"4B", x"42", x"1A", x"5F", x"E1", x"E5", x"66", x"C5", -- 0x5EC8,
      x"2E", x"00", x"55", x"06", x"08", x"29", x"30", x"01", -- 0x5ED0,
      x"19", x"10", x"FA", x"C1", x"EB", x"7B", x"02", x"03", -- 0x5ED8,
      x"7A", x"02", x"C1", x"C5", x"AF", x"02", x"DD", x"7E", -- 0x5EE0,
      x"04", x"DD", x"86", x"08", x"6F", x"DD", x"7E", x"05", -- 0x5EE8,
      x"DD", x"8E", x"09", x"67", x"DD", x"7E", x"06", x"DD", -- 0x5EF0,
      x"8E", x"0A", x"5F", x"DD", x"7E", x"07", x"DD", x"8E", -- 0x5EF8,
      x"0B", x"57", x"DD", x"F9", x"DD", x"E1", x"C9", x"DD", -- 0x5F00,
      x"E5", x"DD", x"21", x"00", x"00", x"DD", x"39", x"3B", -- 0x5F08,
      x"01", x"00", x"00", x"11", x"00", x"00", x"DD", x"36", -- 0x5F10,
      x"FF", x"20", x"DD", x"7E", x"07", x"CB", x"07", x"E6", -- 0x5F18,
      x"01", x"6F", x"DD", x"CB", x"04", x"26", x"DD", x"CB", -- 0x5F20,
      x"05", x"16", x"DD", x"CB", x"06", x"16", x"DD", x"CB", -- 0x5F28,
      x"07", x"16", x"CB", x"21", x"CB", x"10", x"CB", x"13", -- 0x5F30,
      x"CB", x"12", x"CB", x"45", x"28", x"02", x"CB", x"C1", -- 0x5F38,
      x"79", x"DD", x"96", x"08", x"78", x"DD", x"9E", x"09", -- 0x5F40,
      x"7B", x"DD", x"9E", x"0A", x"7A", x"DD", x"9E", x"0B", -- 0x5F48,
      x"38", x"2E", x"79", x"DD", x"96", x"08", x"4F", x"78", -- 0x5F50,
      x"DD", x"9E", x"09", x"47", x"7B", x"DD", x"9E", x"0A", -- 0x5F58,
      x"5F", x"7A", x"DD", x"9E", x"0B", x"57", x"DD", x"7E", -- 0x5F60,
      x"04", x"F6", x"01", x"DD", x"77", x"04", x"DD", x"7E", -- 0x5F68,
      x"05", x"DD", x"77", x"05", x"DD", x"7E", x"06", x"DD", -- 0x5F70,
      x"77", x"06", x"DD", x"7E", x"07", x"DD", x"77", x"07", -- 0x5F78,
      x"DD", x"35", x"FF", x"DD", x"7E", x"FF", x"B7", x"20", -- 0x5F80,
      x"91", x"DD", x"6E", x"04", x"DD", x"66", x"05", x"DD", -- 0x5F88,
      x"5E", x"06", x"DD", x"56", x"07", x"33", x"DD", x"E1", -- 0x5F90,
      x"C9", x"00", x"00", x"20", x"00", x"00", x"00", x"00", -- 0x5F98,
      x"00", x"00", x"00", x"00", x"00", x"BE", x"17", x"DE", -- 0x5FA0,
      x"17", x"CE", x"17", x"00", x"00", x"00", x"00", x"01", -- 0x5FA8,
      x"01", x"17", x"00", x"78", x"B1", x"CA", x"41", x"0C", -- 0x5FB0,
      x"11", x"44", x"73", x"21", x"99", x"5F", x"ED", x"B0", -- 0x5FB8,
      x"FD", x"21", x"C1", x"66", x"FD", x"36", x"00", x"FF", -- 0x5FC0,
      x"FD", x"21", x"C2", x"66", x"FD", x"36", x"00", x"00", -- 0x5FC8,
      x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FD0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FD8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FE0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FE8,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FF0,
      x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", -- 0x5FF8
   );

begin
   process(clock_i)
   begin
      if rising_edge(clock_i) then
         if we_n_i = '1' then
            ram_q(to_integer(unsigned(addr_i))) <= data_i;
         end if;
         data_o <= ram_q(to_integer(unsigned(addr_i)));
      end if;
   end process;

end rtl;
